WIDTH=16;
DEPTH=9;
ADDRESS_RADIX=UNS;
DATA_RADIX=HEX;

CONTENT BEGIN
	0 : fffe;
	1 : 0000;
	2 : 0001;
	3 : 0000;
	4 : 0000;
	5 : 0000;
	6 : 0000;
	7 : 0000;
	8 : 0000;
END;