`timescale 1ns / 1ps
module instruction_rom #( parameter SIZE = 32)
(
	input logic CLK,
	input logic Reset,
	input logic [SIZE-1:0] Address,
	output logic [SIZE-1:0] Instr
);
always@(posedge CLK) begin
	if( Reset ) Instr <= 48'bx;
	else begin
		case (Address/48'd4)
			48'H000000000000: Instr <= 48'He83004000000;
			48'H000000000001: Instr <= 48'He14002000001;
			48'H000000000002: Instr <= 48'He83006000001;
			48'H000000000003: Instr <= 48'He14042000001;
			48'H000000000004: Instr <= 48'He83008000001;
			48'H000000000005: Instr <= 48'He02042000001;
			48'H000000000006: Instr <= 48'He9300a000000;
			48'H000000000007: Instr <= 48'He1f980000280;
			48'H000000000008: Instr <= 48'H0a0780000012;
			48'H000000000009: Instr <= 48'He1f9c00001e0;
			48'H00000000000a: Instr <= 48'H0a0780000013;
			48'H00000000000b: Instr <= 48'He04210000007;
			48'H00000000000c: Instr <= 48'Hec3212000006;
			48'H00000000000d: Instr <= 48'He14210000001;
			48'H00000000000e: Instr <= 48'Hec3214000006;
			48'H00000000000f: Instr <= 48'He14210000001;
			48'H000000000010: Instr <= 48'Hec3216000006;
			48'H000000000011: Instr <= 48'He0c252000002;
			48'H000000000012: Instr <= 48'He0c294000003;
			48'H000000000013: Instr <= 48'He0c2d6000004;
			48'H000000000014: Instr <= 48'He0425200000a;
			48'H000000000015: Instr <= 48'He0425200000b;
			48'H000000000016: Instr <= 48'He0d252000005;
			48'H000000000017: Instr <= 48'Hea4258000000;
			48'H000000000018: Instr <= 48'He02210000008;
			48'H000000000019: Instr <= 48'He1418c000001;
			48'H00000000001a: Instr <= 48'He14318000004;
			48'H00000000001b: Instr <= 48'He403c0ffffea;
			48'H00000000001c: Instr <= 48'He141ce000001;
			48'H00000000001d: Instr <= 48'He0218c000006;
			48'H00000000001e: Instr <= 48'He403c0ffffe7;
			48'H00000000001f: Instr <= 48'He0435a00000d;
			default: Instr <= 48'bx;
		endcase
	end
end
endmodule
