`timescale 1ns / 1ps
module mem_pic #( parameter SIZE = 8 )
(
	input logic CLK,
	input logic [31:0] ADDRESS,
	output logic [SIZE-1:0] READ
);

always_ff@( posedge CLK ) begin
	case( ADDRESS )
		
		32'H00000000: READ <= 8'Hb3;
		32'H00000001: READ <= 8'Hb6;
		32'H00000002: READ <= 8'Hb8;
		32'H00000003: READ <= 8'Hbb;
		32'H00000004: READ <= 8'Hbe;
		32'H00000005: READ <= 8'Hc1;
		32'H00000006: READ <= 8'Hc5;
		32'H00000007: READ <= 8'Hc8;
		32'H00000008: READ <= 8'Hcb;
		32'H00000009: READ <= 8'Hce;
		32'H0000000a: READ <= 8'Hd2;
		32'H0000000b: READ <= 8'Hd5;
		32'H0000000c: READ <= 8'Hd6;
		32'H0000000d: READ <= 8'Hda;
		32'H0000000e: READ <= 8'Hdc;
		32'H0000000f: READ <= 8'Hdf;
		32'H00000010: READ <= 8'He1;
		32'H00000011: READ <= 8'He4;
		32'H00000012: READ <= 8'He6;
		32'H00000013: READ <= 8'He8;
		32'H00000014: READ <= 8'He9;
		32'H00000015: READ <= 8'Hea;
		32'H00000016: READ <= 8'Heb;
		32'H00000017: READ <= 8'Hec;
		32'H00000018: READ <= 8'Hee;
		32'H00000019: READ <= 8'Hee;
		32'H0000001a: READ <= 8'Hef;
		32'H0000001b: READ <= 8'Hef;
		32'H0000001c: READ <= 8'Hf0;
		32'H0000001d: READ <= 8'Hf1;
		32'H0000001e: READ <= 8'Hf2;
		32'H0000001f: READ <= 8'Hf2;
		32'H00000020: READ <= 8'Hf2;
		32'H00000021: READ <= 8'Hf2;
		32'H00000022: READ <= 8'Hf1;
		32'H00000023: READ <= 8'Hf0;
		32'H00000024: READ <= 8'Hef;
		32'H00000025: READ <= 8'Hee;
		32'H00000026: READ <= 8'Hed;
		32'H00000027: READ <= 8'Hea;
		32'H00000028: READ <= 8'He9;
		32'H00000029: READ <= 8'He8;
		32'H0000002a: READ <= 8'He6;
		32'H0000002b: READ <= 8'He2;
		32'H0000002c: READ <= 8'He0;
		32'H0000002d: READ <= 8'Hdc;
		32'H0000002e: READ <= 8'Hd7;
		32'H0000002f: READ <= 8'Hd3;
		32'H00000030: READ <= 8'Hce;
		32'H00000031: READ <= 8'Hc9;
		32'H00000032: READ <= 8'Hc3;
		32'H00000033: READ <= 8'Hbc;
		32'H00000034: READ <= 8'Hb3;
		32'H00000035: READ <= 8'Hac;
		32'H00000036: READ <= 8'Ha6;
		32'H00000037: READ <= 8'Ha1;
		32'H00000038: READ <= 8'H9f;
		32'H00000039: READ <= 8'H9d;
		32'H0000003a: READ <= 8'H9c;
		32'H0000003b: READ <= 8'H9b;
		32'H0000003c: READ <= 8'H9b;
		32'H0000003d: READ <= 8'H9b;
		32'H0000003e: READ <= 8'H9a;
		32'H0000003f: READ <= 8'H9b;
		32'H00000040: READ <= 8'H9b;
		32'H00000041: READ <= 8'H9b;
		32'H00000042: READ <= 8'H9c;
		32'H00000043: READ <= 8'H9d;
		32'H00000044: READ <= 8'H9d;
		32'H00000045: READ <= 8'H9d;
		32'H00000046: READ <= 8'H9d;
		32'H00000047: READ <= 8'H9d;
		32'H00000048: READ <= 8'H9e;
		32'H00000049: READ <= 8'H9d;
		32'H0000004a: READ <= 8'H9e;
		32'H0000004b: READ <= 8'H9f;
		32'H0000004c: READ <= 8'H9f;
		32'H0000004d: READ <= 8'H9f;
		32'H0000004e: READ <= 8'Ha0;
		32'H0000004f: READ <= 8'Ha1;
		32'H00000050: READ <= 8'Ha1;
		32'H00000051: READ <= 8'Ha2;
		32'H00000052: READ <= 8'Ha2;
		32'H00000053: READ <= 8'Ha3;
		32'H00000054: READ <= 8'Ha3;
		32'H00000055: READ <= 8'Ha3;
		32'H00000056: READ <= 8'Ha4;
		32'H00000057: READ <= 8'Ha4;
		32'H00000058: READ <= 8'Ha4;
		32'H00000059: READ <= 8'Ha4;
		32'H0000005a: READ <= 8'Ha4;
		32'H0000005b: READ <= 8'Ha3;
		32'H0000005c: READ <= 8'Ha4;
		32'H0000005d: READ <= 8'Ha4;
		32'H0000005e: READ <= 8'Ha5;
		32'H0000005f: READ <= 8'Ha5;
		32'H00000060: READ <= 8'Ha6;
		32'H00000061: READ <= 8'Ha7;
		32'H00000062: READ <= 8'Ha7;
		32'H00000063: READ <= 8'Ha8;
		
		32'H00010000: READ <= 8'Hb3;
		32'H00010001: READ <= 8'Hb5;
		32'H00010002: READ <= 8'Hb7;
		32'H00010003: READ <= 8'Hb9;
		32'H00010004: READ <= 8'Hbc;
		32'H00010005: READ <= 8'Hbf;
		32'H00010006: READ <= 8'Hc3;
		32'H00010007: READ <= 8'Hc6;
		32'H00010008: READ <= 8'Hc9;
		32'H00010009: READ <= 8'Hcd;
		32'H0001000a: READ <= 8'Hd1;
		32'H0001000b: READ <= 8'Hd3;
		32'H0001000c: READ <= 8'Hd6;
		32'H0001000d: READ <= 8'Hd9;
		32'H0001000e: READ <= 8'Hdb;
		32'H0001000f: READ <= 8'Hde;
		32'H00010010: READ <= 8'He0;
		32'H00010011: READ <= 8'He4;
		32'H00010012: READ <= 8'He6;
		32'H00010013: READ <= 8'He8;
		32'H00010014: READ <= 8'He9;
		32'H00010015: READ <= 8'Hea;
		32'H00010016: READ <= 8'Hec;
		32'H00010017: READ <= 8'Hec;
		32'H00010018: READ <= 8'Hee;
		32'H00010019: READ <= 8'Hee;
		32'H0001001a: READ <= 8'Hef;
		32'H0001001b: READ <= 8'Hf0;
		32'H0001001c: READ <= 8'Hf0;
		32'H0001001d: READ <= 8'Hf2;
		32'H0001001e: READ <= 8'Hf2;
		32'H0001001f: READ <= 8'Hf2;
		32'H00010020: READ <= 8'Hf2;
		32'H00010021: READ <= 8'Hf2;
		32'H00010022: READ <= 8'Hf2;
		32'H00010023: READ <= 8'Hf0;
		32'H00010024: READ <= 8'Hef;
		32'H00010025: READ <= 8'Hee;
		32'H00010026: READ <= 8'Hec;
		32'H00010027: READ <= 8'Heb;
		32'H00010028: READ <= 8'He9;
		32'H00010029: READ <= 8'He9;
		32'H0001002a: READ <= 8'He7;
		32'H0001002b: READ <= 8'He3;
		32'H0001002c: READ <= 8'He0;
		32'H0001002d: READ <= 8'Hdc;
		32'H0001002e: READ <= 8'Hd8;
		32'H0001002f: READ <= 8'Hd4;
		32'H00010030: READ <= 8'Hd0;
		32'H00010031: READ <= 8'Hcb;
		32'H00010032: READ <= 8'Hc5;
		32'H00010033: READ <= 8'Hbd;
		32'H00010034: READ <= 8'Hb4;
		32'H00010035: READ <= 8'Had;
		32'H00010036: READ <= 8'Ha6;
		32'H00010037: READ <= 8'Ha1;
		32'H00010038: READ <= 8'H9e;
		32'H00010039: READ <= 8'H9c;
		32'H0001003a: READ <= 8'H9b;
		32'H0001003b: READ <= 8'H9a;
		32'H0001003c: READ <= 8'H9b;
		32'H0001003d: READ <= 8'H9a;
		32'H0001003e: READ <= 8'H99;
		32'H0001003f: READ <= 8'H99;
		32'H00010040: READ <= 8'H9a;
		32'H00010041: READ <= 8'H9b;
		32'H00010042: READ <= 8'H9a;
		32'H00010043: READ <= 8'H9b;
		32'H00010044: READ <= 8'H9c;
		32'H00010045: READ <= 8'H9c;
		32'H00010046: READ <= 8'H9d;
		32'H00010047: READ <= 8'H9c;
		32'H00010048: READ <= 8'H9c;
		32'H00010049: READ <= 8'H9c;
		32'H0001004a: READ <= 8'H9c;
		32'H0001004b: READ <= 8'H9d;
		32'H0001004c: READ <= 8'H9e;
		32'H0001004d: READ <= 8'H9e;
		32'H0001004e: READ <= 8'Ha0;
		32'H0001004f: READ <= 8'Ha0;
		32'H00010050: READ <= 8'Ha0;
		32'H00010051: READ <= 8'Ha1;
		32'H00010052: READ <= 8'Ha1;
		32'H00010053: READ <= 8'Ha2;
		32'H00010054: READ <= 8'Ha3;
		32'H00010055: READ <= 8'Ha3;
		32'H00010056: READ <= 8'Ha2;
		32'H00010057: READ <= 8'Ha3;
		32'H00010058: READ <= 8'Ha3;
		32'H00010059: READ <= 8'Ha3;
		32'H0001005a: READ <= 8'Ha3;
		32'H0001005b: READ <= 8'Ha3;
		32'H0001005c: READ <= 8'Ha3;
		32'H0001005d: READ <= 8'Ha3;
		32'H0001005e: READ <= 8'Ha4;
		32'H0001005f: READ <= 8'Ha4;
		32'H00010060: READ <= 8'Ha6;
		32'H00010061: READ <= 8'Ha6;
		32'H00010062: READ <= 8'Ha6;
		32'H00010063: READ <= 8'Ha6;
		
		32'H00020000: READ <= 8'Hb1;
		32'H00020001: READ <= 8'Hb3;
		32'H00020002: READ <= 8'Hb6;
		32'H00020003: READ <= 8'Hb8;
		32'H00020004: READ <= 8'Hba;
		32'H00020005: READ <= 8'Hbd;
		32'H00020006: READ <= 8'Hc1;
		32'H00020007: READ <= 8'Hc5;
		32'H00020008: READ <= 8'Hc8;
		32'H00020009: READ <= 8'Hcc;
		32'H0002000a: READ <= 8'Hcf;
		32'H0002000b: READ <= 8'Hd2;
		32'H0002000c: READ <= 8'Hd5;
		32'H0002000d: READ <= 8'Hd8;
		32'H0002000e: READ <= 8'Hda;
		32'H0002000f: READ <= 8'Hdd;
		32'H00020010: READ <= 8'He0;
		32'H00020011: READ <= 8'He3;
		32'H00020012: READ <= 8'He5;
		32'H00020013: READ <= 8'He7;
		32'H00020014: READ <= 8'He9;
		32'H00020015: READ <= 8'Hea;
		32'H00020016: READ <= 8'Heb;
		32'H00020017: READ <= 8'Hec;
		32'H00020018: READ <= 8'Hee;
		32'H00020019: READ <= 8'Hee;
		32'H0002001a: READ <= 8'Hef;
		32'H0002001b: READ <= 8'Hef;
		32'H0002001c: READ <= 8'Hf1;
		32'H0002001d: READ <= 8'Hf2;
		32'H0002001e: READ <= 8'Hf2;
		32'H0002001f: READ <= 8'Hf2;
		32'H00020020: READ <= 8'Hf2;
		32'H00020021: READ <= 8'Hf2;
		32'H00020022: READ <= 8'Hf2;
		32'H00020023: READ <= 8'Hf1;
		32'H00020024: READ <= 8'Hef;
		32'H00020025: READ <= 8'Hee;
		32'H00020026: READ <= 8'Hed;
		32'H00020027: READ <= 8'Hec;
		32'H00020028: READ <= 8'Hea;
		32'H00020029: READ <= 8'Heb;
		32'H0002002a: READ <= 8'Hea;
		32'H0002002b: READ <= 8'He6;
		32'H0002002c: READ <= 8'He1;
		32'H0002002d: READ <= 8'Hdd;
		32'H0002002e: READ <= 8'Hda;
		32'H0002002f: READ <= 8'Hd5;
		32'H00020030: READ <= 8'Hd1;
		32'H00020031: READ <= 8'Hcc;
		32'H00020032: READ <= 8'Hc6;
		32'H00020033: READ <= 8'Hbe;
		32'H00020034: READ <= 8'Hb6;
		32'H00020035: READ <= 8'Had;
		32'H00020036: READ <= 8'Ha7;
		32'H00020037: READ <= 8'Ha1;
		32'H00020038: READ <= 8'H9e;
		32'H00020039: READ <= 8'H9c;
		32'H0002003a: READ <= 8'H9a;
		32'H0002003b: READ <= 8'H9a;
		32'H0002003c: READ <= 8'H98;
		32'H0002003d: READ <= 8'H98;
		32'H0002003e: READ <= 8'H98;
		32'H0002003f: READ <= 8'H98;
		32'H00020040: READ <= 8'H99;
		32'H00020041: READ <= 8'H99;
		32'H00020042: READ <= 8'H99;
		32'H00020043: READ <= 8'H9a;
		32'H00020044: READ <= 8'H9a;
		32'H00020045: READ <= 8'H9b;
		32'H00020046: READ <= 8'H9b;
		32'H00020047: READ <= 8'H9b;
		32'H00020048: READ <= 8'H9a;
		32'H00020049: READ <= 8'H9b;
		32'H0002004a: READ <= 8'H9b;
		32'H0002004b: READ <= 8'H9c;
		32'H0002004c: READ <= 8'H9d;
		32'H0002004d: READ <= 8'H9d;
		32'H0002004e: READ <= 8'H9e;
		32'H0002004f: READ <= 8'H9e;
		32'H00020050: READ <= 8'H9f;
		32'H00020051: READ <= 8'H9f;
		32'H00020052: READ <= 8'Ha0;
		32'H00020053: READ <= 8'Ha1;
		32'H00020054: READ <= 8'Ha2;
		32'H00020055: READ <= 8'Ha1;
		32'H00020056: READ <= 8'Ha1;
		32'H00020057: READ <= 8'Ha2;
		32'H00020058: READ <= 8'Ha1;
		32'H00020059: READ <= 8'Ha2;
		32'H0002005a: READ <= 8'Ha2;
		32'H0002005b: READ <= 8'Ha1;
		32'H0002005c: READ <= 8'Ha2;
		32'H0002005d: READ <= 8'Ha3;
		32'H0002005e: READ <= 8'Ha3;
		32'H0002005f: READ <= 8'Ha3;
		32'H00020060: READ <= 8'Ha4;
		32'H00020061: READ <= 8'Ha5;
		32'H00020062: READ <= 8'Ha5;
		32'H00020063: READ <= 8'Ha6;
		
		32'H00030000: READ <= 8'Haf;
		32'H00030001: READ <= 8'Hb3;
		32'H00030002: READ <= 8'Hb5;
		32'H00030003: READ <= 8'Hb6;
		32'H00030004: READ <= 8'Hb9;
		32'H00030005: READ <= 8'Hbb;
		32'H00030006: READ <= 8'Hbf;
		32'H00030007: READ <= 8'Hc3;
		32'H00030008: READ <= 8'Hc6;
		32'H00030009: READ <= 8'Hca;
		32'H0003000a: READ <= 8'Hcd;
		32'H0003000b: READ <= 8'Hd1;
		32'H0003000c: READ <= 8'Hd3;
		32'H0003000d: READ <= 8'Hd6;
		32'H0003000e: READ <= 8'Hda;
		32'H0003000f: READ <= 8'Hdc;
		32'H00030010: READ <= 8'Hdf;
		32'H00030011: READ <= 8'He2;
		32'H00030012: READ <= 8'He5;
		32'H00030013: READ <= 8'He7;
		32'H00030014: READ <= 8'He8;
		32'H00030015: READ <= 8'Hea;
		32'H00030016: READ <= 8'Heb;
		32'H00030017: READ <= 8'Heb;
		32'H00030018: READ <= 8'Hed;
		32'H00030019: READ <= 8'Hee;
		32'H0003001a: READ <= 8'Hee;
		32'H0003001b: READ <= 8'Hf0;
		32'H0003001c: READ <= 8'Hf1;
		32'H0003001d: READ <= 8'Hf2;
		32'H0003001e: READ <= 8'Hf2;
		32'H0003001f: READ <= 8'Hf3;
		32'H00030020: READ <= 8'Hf3;
		32'H00030021: READ <= 8'Hf2;
		32'H00030022: READ <= 8'Hf2;
		32'H00030023: READ <= 8'Hf1;
		32'H00030024: READ <= 8'Hef;
		32'H00030025: READ <= 8'Hee;
		32'H00030026: READ <= 8'Hed;
		32'H00030027: READ <= 8'Hed;
		32'H00030028: READ <= 8'Hed;
		32'H00030029: READ <= 8'Hee;
		32'H0003002a: READ <= 8'Hee;
		32'H0003002b: READ <= 8'Hec;
		32'H0003002c: READ <= 8'He3;
		32'H0003002d: READ <= 8'Hde;
		32'H0003002e: READ <= 8'Hdb;
		32'H0003002f: READ <= 8'Hd7;
		32'H00030030: READ <= 8'Hd1;
		32'H00030031: READ <= 8'Hcd;
		32'H00030032: READ <= 8'Hc7;
		32'H00030033: READ <= 8'Hc0;
		32'H00030034: READ <= 8'Hb7;
		32'H00030035: READ <= 8'Haf;
		32'H00030036: READ <= 8'Ha7;
		32'H00030037: READ <= 8'Ha2;
		32'H00030038: READ <= 8'H9e;
		32'H00030039: READ <= 8'H9b;
		32'H0003003a: READ <= 8'H9a;
		32'H0003003b: READ <= 8'H99;
		32'H0003003c: READ <= 8'H97;
		32'H0003003d: READ <= 8'H96;
		32'H0003003e: READ <= 8'H97;
		32'H0003003f: READ <= 8'H97;
		32'H00030040: READ <= 8'H97;
		32'H00030041: READ <= 8'H98;
		32'H00030042: READ <= 8'H98;
		32'H00030043: READ <= 8'H99;
		32'H00030044: READ <= 8'H99;
		32'H00030045: READ <= 8'H9a;
		32'H00030046: READ <= 8'H9a;
		32'H00030047: READ <= 8'H9a;
		32'H00030048: READ <= 8'H99;
		32'H00030049: READ <= 8'H9a;
		32'H0003004a: READ <= 8'H9a;
		32'H0003004b: READ <= 8'H9b;
		32'H0003004c: READ <= 8'H9b;
		32'H0003004d: READ <= 8'H9c;
		32'H0003004e: READ <= 8'H9d;
		32'H0003004f: READ <= 8'H9e;
		32'H00030050: READ <= 8'H9e;
		32'H00030051: READ <= 8'H9f;
		32'H00030052: READ <= 8'H9f;
		32'H00030053: READ <= 8'Ha0;
		32'H00030054: READ <= 8'Ha0;
		32'H00030055: READ <= 8'Ha0;
		32'H00030056: READ <= 8'Ha0;
		32'H00030057: READ <= 8'Ha1;
		32'H00030058: READ <= 8'Ha1;
		32'H00030059: READ <= 8'Ha1;
		32'H0003005a: READ <= 8'Ha1;
		32'H0003005b: READ <= 8'Ha1;
		32'H0003005c: READ <= 8'Ha1;
		32'H0003005d: READ <= 8'Ha1;
		32'H0003005e: READ <= 8'Ha1;
		32'H0003005f: READ <= 8'Ha2;
		32'H00030060: READ <= 8'Ha3;
		32'H00030061: READ <= 8'Ha4;
		32'H00030062: READ <= 8'Ha4;
		32'H00030063: READ <= 8'Ha5;
		
		32'H00040000: READ <= 8'Had;
		32'H00040001: READ <= 8'Hb1;
		32'H00040002: READ <= 8'Hb3;
		32'H00040003: READ <= 8'Hb4;
		32'H00040004: READ <= 8'Hb6;
		32'H00040005: READ <= 8'Hba;
		32'H00040006: READ <= 8'Hbe;
		32'H00040007: READ <= 8'Hc1;
		32'H00040008: READ <= 8'Hc4;
		32'H00040009: READ <= 8'Hc8;
		32'H0004000a: READ <= 8'Hcc;
		32'H0004000b: READ <= 8'Hd0;
		32'H0004000c: READ <= 8'Hd2;
		32'H0004000d: READ <= 8'Hd5;
		32'H0004000e: READ <= 8'Hd8;
		32'H0004000f: READ <= 8'Hdc;
		32'H00040010: READ <= 8'Hdf;
		32'H00040011: READ <= 8'He1;
		32'H00040012: READ <= 8'He4;
		32'H00040013: READ <= 8'He7;
		32'H00040014: READ <= 8'He8;
		32'H00040015: READ <= 8'He9;
		32'H00040016: READ <= 8'Heb;
		32'H00040017: READ <= 8'Hec;
		32'H00040018: READ <= 8'Hed;
		32'H00040019: READ <= 8'Hee;
		32'H0004001a: READ <= 8'Hef;
		32'H0004001b: READ <= 8'Hf0;
		32'H0004001c: READ <= 8'Hf1;
		32'H0004001d: READ <= 8'Hf2;
		32'H0004001e: READ <= 8'Hf2;
		32'H0004001f: READ <= 8'Hf2;
		32'H00040020: READ <= 8'Hf3;
		32'H00040021: READ <= 8'Hf2;
		32'H00040022: READ <= 8'Hf2;
		32'H00040023: READ <= 8'Hf1;
		32'H00040024: READ <= 8'Hf0;
		32'H00040025: READ <= 8'Hf0;
		32'H00040026: READ <= 8'Hf0;
		32'H00040027: READ <= 8'Hef;
		32'H00040028: READ <= 8'Heb;
		32'H00040029: READ <= 8'He4;
		32'H0004002a: READ <= 8'Hdc;
		32'H0004002b: READ <= 8'Hdf;
		32'H0004002c: READ <= 8'He2;
		32'H0004002d: READ <= 8'He4;
		32'H0004002e: READ <= 8'He1;
		32'H0004002f: READ <= 8'Hde;
		32'H00040030: READ <= 8'Hda;
		32'H00040031: READ <= 8'Hd1;
		32'H00040032: READ <= 8'Hcc;
		32'H00040033: READ <= 8'Hc2;
		32'H00040034: READ <= 8'Hb9;
		32'H00040035: READ <= 8'Haf;
		32'H00040036: READ <= 8'Ha8;
		32'H00040037: READ <= 8'Ha2;
		32'H00040038: READ <= 8'H9e;
		32'H00040039: READ <= 8'H9a;
		32'H0004003a: READ <= 8'H99;
		32'H0004003b: READ <= 8'H98;
		32'H0004003c: READ <= 8'H98;
		32'H0004003d: READ <= 8'H96;
		32'H0004003e: READ <= 8'H96;
		32'H0004003f: READ <= 8'H96;
		32'H00040040: READ <= 8'H95;
		32'H00040041: READ <= 8'H96;
		32'H00040042: READ <= 8'H97;
		32'H00040043: READ <= 8'H97;
		32'H00040044: READ <= 8'H98;
		32'H00040045: READ <= 8'H99;
		32'H00040046: READ <= 8'H99;
		32'H00040047: READ <= 8'H99;
		32'H00040048: READ <= 8'H99;
		32'H00040049: READ <= 8'H99;
		32'H0004004a: READ <= 8'H99;
		32'H0004004b: READ <= 8'H9a;
		32'H0004004c: READ <= 8'H99;
		32'H0004004d: READ <= 8'H9b;
		32'H0004004e: READ <= 8'H9c;
		32'H0004004f: READ <= 8'H9c;
		32'H00040050: READ <= 8'H9d;
		32'H00040051: READ <= 8'H9e;
		32'H00040052: READ <= 8'H9d;
		32'H00040053: READ <= 8'H9e;
		32'H00040054: READ <= 8'H9e;
		32'H00040055: READ <= 8'H9f;
		32'H00040056: READ <= 8'H9f;
		32'H00040057: READ <= 8'H9f;
		32'H00040058: READ <= 8'Ha0;
		32'H00040059: READ <= 8'Ha0;
		32'H0004005a: READ <= 8'Ha0;
		32'H0004005b: READ <= 8'Ha1;
		32'H0004005c: READ <= 8'Ha0;
		32'H0004005d: READ <= 8'Ha0;
		32'H0004005e: READ <= 8'Ha1;
		32'H0004005f: READ <= 8'Ha2;
		32'H00040060: READ <= 8'Ha2;
		32'H00040061: READ <= 8'Ha2;
		32'H00040062: READ <= 8'Ha3;
		32'H00040063: READ <= 8'Ha4;
		
		32'H00050000: READ <= 8'Hab;
		32'H00050001: READ <= 8'Haf;
		32'H00050002: READ <= 8'Hb1;
		32'H00050003: READ <= 8'Hb3;
		32'H00050004: READ <= 8'Hb5;
		32'H00050005: READ <= 8'Hb8;
		32'H00050006: READ <= 8'Hbb;
		32'H00050007: READ <= 8'Hbf;
		32'H00050008: READ <= 8'Hc2;
		32'H00050009: READ <= 8'Hc6;
		32'H0005000a: READ <= 8'Hcb;
		32'H0005000b: READ <= 8'Hce;
		32'H0005000c: READ <= 8'Hd2;
		32'H0005000d: READ <= 8'Hd4;
		32'H0005000e: READ <= 8'Hd7;
		32'H0005000f: READ <= 8'Hdb;
		32'H00050010: READ <= 8'Hde;
		32'H00050011: READ <= 8'He1;
		32'H00050012: READ <= 8'He4;
		32'H00050013: READ <= 8'He6;
		32'H00050014: READ <= 8'He8;
		32'H00050015: READ <= 8'He9;
		32'H00050016: READ <= 8'Heb;
		32'H00050017: READ <= 8'Hec;
		32'H00050018: READ <= 8'Hed;
		32'H00050019: READ <= 8'Hee;
		32'H0005001a: READ <= 8'Hef;
		32'H0005001b: READ <= 8'Hf1;
		32'H0005001c: READ <= 8'Hf1;
		32'H0005001d: READ <= 8'Hf2;
		32'H0005001e: READ <= 8'Hf3;
		32'H0005001f: READ <= 8'Hf3;
		32'H00050020: READ <= 8'Hf3;
		32'H00050021: READ <= 8'Hf2;
		32'H00050022: READ <= 8'Hf3;
		32'H00050023: READ <= 8'Hf1;
		32'H00050024: READ <= 8'Hf4;
		32'H00050025: READ <= 8'Hef;
		32'H00050026: READ <= 8'Hd5;
		32'H00050027: READ <= 8'Hca;
		32'H00050028: READ <= 8'Hc2;
		32'H00050029: READ <= 8'Hc2;
		32'H0005002a: READ <= 8'Hbd;
		32'H0005002b: READ <= 8'Hb6;
		32'H0005002c: READ <= 8'Hbc;
		32'H0005002d: READ <= 8'Hc6;
		32'H0005002e: READ <= 8'Hcc;
		32'H0005002f: READ <= 8'Hbc;
		32'H00050030: READ <= 8'Hc1;
		32'H00050031: READ <= 8'Hc8;
		32'H00050032: READ <= 8'Hba;
		32'H00050033: READ <= 8'Hc2;
		32'H00050034: READ <= 8'Hb8;
		32'H00050035: READ <= 8'Hb1;
		32'H00050036: READ <= 8'Ha9;
		32'H00050037: READ <= 8'Ha2;
		32'H00050038: READ <= 8'H9d;
		32'H00050039: READ <= 8'H9a;
		32'H0005003a: READ <= 8'H98;
		32'H0005003b: READ <= 8'H97;
		32'H0005003c: READ <= 8'H97;
		32'H0005003d: READ <= 8'H95;
		32'H0005003e: READ <= 8'H95;
		32'H0005003f: READ <= 8'H95;
		32'H00050040: READ <= 8'H95;
		32'H00050041: READ <= 8'H96;
		32'H00050042: READ <= 8'H96;
		32'H00050043: READ <= 8'H96;
		32'H00050044: READ <= 8'H97;
		32'H00050045: READ <= 8'H98;
		32'H00050046: READ <= 8'H97;
		32'H00050047: READ <= 8'H97;
		32'H00050048: READ <= 8'H97;
		32'H00050049: READ <= 8'H98;
		32'H0005004a: READ <= 8'H98;
		32'H0005004b: READ <= 8'H99;
		32'H0005004c: READ <= 8'H99;
		32'H0005004d: READ <= 8'H9a;
		32'H0005004e: READ <= 8'H9b;
		32'H0005004f: READ <= 8'H9c;
		32'H00050050: READ <= 8'H9c;
		32'H00050051: READ <= 8'H9d;
		32'H00050052: READ <= 8'H9d;
		32'H00050053: READ <= 8'H9d;
		32'H00050054: READ <= 8'H9d;
		32'H00050055: READ <= 8'H9e;
		32'H00050056: READ <= 8'H9e;
		32'H00050057: READ <= 8'H9e;
		32'H00050058: READ <= 8'H9f;
		32'H00050059: READ <= 8'H9f;
		32'H0005005a: READ <= 8'H9f;
		32'H0005005b: READ <= 8'Ha0;
		32'H0005005c: READ <= 8'Ha0;
		32'H0005005d: READ <= 8'Ha0;
		32'H0005005e: READ <= 8'Ha0;
		32'H0005005f: READ <= 8'Ha0;
		32'H00050060: READ <= 8'Ha1;
		32'H00050061: READ <= 8'Ha2;
		32'H00050062: READ <= 8'Ha2;
		32'H00050063: READ <= 8'Ha2;
		
		32'H00060000: READ <= 8'Ha9;
		32'H00060001: READ <= 8'Hac;
		32'H00060002: READ <= 8'Haf;
		32'H00060003: READ <= 8'Hb2;
		32'H00060004: READ <= 8'Hb4;
		32'H00060005: READ <= 8'Hb7;
		32'H00060006: READ <= 8'Hba;
		32'H00060007: READ <= 8'Hbd;
		32'H00060008: READ <= 8'Hc1;
		32'H00060009: READ <= 8'Hc4;
		32'H0006000a: READ <= 8'Hc9;
		32'H0006000b: READ <= 8'Hcd;
		32'H0006000c: READ <= 8'Hd1;
		32'H0006000d: READ <= 8'Hd3;
		32'H0006000e: READ <= 8'Hd6;
		32'H0006000f: READ <= 8'Hd9;
		32'H00060010: READ <= 8'Hdd;
		32'H00060011: READ <= 8'He0;
		32'H00060012: READ <= 8'He3;
		32'H00060013: READ <= 8'He5;
		32'H00060014: READ <= 8'He7;
		32'H00060015: READ <= 8'He9;
		32'H00060016: READ <= 8'Heb;
		32'H00060017: READ <= 8'Hec;
		32'H00060018: READ <= 8'Hed;
		32'H00060019: READ <= 8'Hee;
		32'H0006001a: READ <= 8'Hef;
		32'H0006001b: READ <= 8'Hf0;
		32'H0006001c: READ <= 8'Hf1;
		32'H0006001d: READ <= 8'Hf2;
		32'H0006001e: READ <= 8'Hf3;
		32'H0006001f: READ <= 8'Hf3;
		32'H00060020: READ <= 8'Hf3;
		32'H00060021: READ <= 8'Hf3;
		32'H00060022: READ <= 8'Hf1;
		32'H00060023: READ <= 8'Hf8;
		32'H00060024: READ <= 8'He5;
		32'H00060025: READ <= 8'Hbb;
		32'H00060026: READ <= 8'H9e;
		32'H00060027: READ <= 8'Haa;
		32'H00060028: READ <= 8'Hb3;
		32'H00060029: READ <= 8'Ha8;
		32'H0006002a: READ <= 8'Had;
		32'H0006002b: READ <= 8'Hac;
		32'H0006002c: READ <= 8'H9e;
		32'H0006002d: READ <= 8'Ha3;
		32'H0006002e: READ <= 8'H9b;
		32'H0006002f: READ <= 8'H9e;
		32'H00060030: READ <= 8'H93;
		32'H00060031: READ <= 8'Ha7;
		32'H00060032: READ <= 8'Ha1;
		32'H00060033: READ <= 8'H9e;
		32'H00060034: READ <= 8'Hac;
		32'H00060035: READ <= 8'Hb6;
		32'H00060036: READ <= 8'Hac;
		32'H00060037: READ <= 8'Ha2;
		32'H00060038: READ <= 8'H9d;
		32'H00060039: READ <= 8'H99;
		32'H0006003a: READ <= 8'H98;
		32'H0006003b: READ <= 8'H96;
		32'H0006003c: READ <= 8'H96;
		32'H0006003d: READ <= 8'H95;
		32'H0006003e: READ <= 8'H94;
		32'H0006003f: READ <= 8'H94;
		32'H00060040: READ <= 8'H93;
		32'H00060041: READ <= 8'H94;
		32'H00060042: READ <= 8'H95;
		32'H00060043: READ <= 8'H95;
		32'H00060044: READ <= 8'H96;
		32'H00060045: READ <= 8'H96;
		32'H00060046: READ <= 8'H96;
		32'H00060047: READ <= 8'H96;
		32'H00060048: READ <= 8'H96;
		32'H00060049: READ <= 8'H97;
		32'H0006004a: READ <= 8'H97;
		32'H0006004b: READ <= 8'H97;
		32'H0006004c: READ <= 8'H99;
		32'H0006004d: READ <= 8'H99;
		32'H0006004e: READ <= 8'H9a;
		32'H0006004f: READ <= 8'H9b;
		32'H00060050: READ <= 8'H9b;
		32'H00060051: READ <= 8'H9b;
		32'H00060052: READ <= 8'H9c;
		32'H00060053: READ <= 8'H9c;
		32'H00060054: READ <= 8'H9c;
		32'H00060055: READ <= 8'H9e;
		32'H00060056: READ <= 8'H9e;
		32'H00060057: READ <= 8'H9e;
		32'H00060058: READ <= 8'H9e;
		32'H00060059: READ <= 8'H9e;
		32'H0006005a: READ <= 8'H9f;
		32'H0006005b: READ <= 8'H9f;
		32'H0006005c: READ <= 8'H9e;
		32'H0006005d: READ <= 8'H9e;
		32'H0006005e: READ <= 8'H9f;
		32'H0006005f: READ <= 8'H9f;
		32'H00060060: READ <= 8'Ha0;
		32'H00060061: READ <= 8'Ha1;
		32'H00060062: READ <= 8'Ha1;
		32'H00060063: READ <= 8'Ha1;
		
		32'H00070000: READ <= 8'Ha7;
		32'H00070001: READ <= 8'Ha9;
		32'H00070002: READ <= 8'Had;
		32'H00070003: READ <= 8'Hb0;
		32'H00070004: READ <= 8'Hb2;
		32'H00070005: READ <= 8'Hb6;
		32'H00070006: READ <= 8'Hb8;
		32'H00070007: READ <= 8'Hbc;
		32'H00070008: READ <= 8'Hc0;
		32'H00070009: READ <= 8'Hc2;
		32'H0007000a: READ <= 8'Hc7;
		32'H0007000b: READ <= 8'Hcc;
		32'H0007000c: READ <= 8'Hd0;
		32'H0007000d: READ <= 8'Hd2;
		32'H0007000e: READ <= 8'Hd5;
		32'H0007000f: READ <= 8'Hd8;
		32'H00070010: READ <= 8'Hdc;
		32'H00070011: READ <= 8'Hdf;
		32'H00070012: READ <= 8'He2;
		32'H00070013: READ <= 8'He5;
		32'H00070014: READ <= 8'He7;
		32'H00070015: READ <= 8'He8;
		32'H00070016: READ <= 8'Hea;
		32'H00070017: READ <= 8'Heb;
		32'H00070018: READ <= 8'Hed;
		32'H00070019: READ <= 8'Hee;
		32'H0007001a: READ <= 8'Hef;
		32'H0007001b: READ <= 8'Hf0;
		32'H0007001c: READ <= 8'Hf1;
		32'H0007001d: READ <= 8'Hf2;
		32'H0007001e: READ <= 8'Hf2;
		32'H0007001f: READ <= 8'Hf3;
		32'H00070020: READ <= 8'Hf3;
		32'H00070021: READ <= 8'Hf5;
		32'H00070022: READ <= 8'Hf7;
		32'H00070023: READ <= 8'Hc8;
		32'H00070024: READ <= 8'Ha8;
		32'H00070025: READ <= 8'Haa;
		32'H00070026: READ <= 8'Ha1;
		32'H00070027: READ <= 8'H88;
		32'H00070028: READ <= 8'Hae;
		32'H00070029: READ <= 8'Ha6;
		32'H0007002a: READ <= 8'Hac;
		32'H0007002b: READ <= 8'Ha3;
		32'H0007002c: READ <= 8'H99;
		32'H0007002d: READ <= 8'H93;
		32'H0007002e: READ <= 8'H91;
		32'H0007002f: READ <= 8'H93;
		32'H00070030: READ <= 8'H82;
		32'H00070031: READ <= 8'H92;
		32'H00070032: READ <= 8'H85;
		32'H00070033: READ <= 8'H77;
		32'H00070034: READ <= 8'H83;
		32'H00070035: READ <= 8'H9b;
		32'H00070036: READ <= 8'Hb2;
		32'H00070037: READ <= 8'Ha7;
		32'H00070038: READ <= 8'H9d;
		32'H00070039: READ <= 8'H9a;
		32'H0007003a: READ <= 8'H97;
		32'H0007003b: READ <= 8'H96;
		32'H0007003c: READ <= 8'H95;
		32'H0007003d: READ <= 8'H94;
		32'H0007003e: READ <= 8'H93;
		32'H0007003f: READ <= 8'H92;
		32'H00070040: READ <= 8'H93;
		32'H00070041: READ <= 8'H93;
		32'H00070042: READ <= 8'H94;
		32'H00070043: READ <= 8'H94;
		32'H00070044: READ <= 8'H94;
		32'H00070045: READ <= 8'H95;
		32'H00070046: READ <= 8'H95;
		32'H00070047: READ <= 8'H95;
		32'H00070048: READ <= 8'H95;
		32'H00070049: READ <= 8'H96;
		32'H0007004a: READ <= 8'H97;
		32'H0007004b: READ <= 8'H97;
		32'H0007004c: READ <= 8'H96;
		32'H0007004d: READ <= 8'H98;
		32'H0007004e: READ <= 8'H99;
		32'H0007004f: READ <= 8'H9a;
		32'H00070050: READ <= 8'H9a;
		32'H00070051: READ <= 8'H9b;
		32'H00070052: READ <= 8'H9b;
		32'H00070053: READ <= 8'H9c;
		32'H00070054: READ <= 8'H9d;
		32'H00070055: READ <= 8'H9d;
		32'H00070056: READ <= 8'H9d;
		32'H00070057: READ <= 8'H9d;
		32'H00070058: READ <= 8'H9d;
		32'H00070059: READ <= 8'H9d;
		32'H0007005a: READ <= 8'H9e;
		32'H0007005b: READ <= 8'H9e;
		32'H0007005c: READ <= 8'H9e;
		32'H0007005d: READ <= 8'H9e;
		32'H0007005e: READ <= 8'H9d;
		32'H0007005f: READ <= 8'H9e;
		32'H00070060: READ <= 8'H9e;
		32'H00070061: READ <= 8'H9f;
		32'H00070062: READ <= 8'Ha0;
		32'H00070063: READ <= 8'Ha0;
		
		32'H00080000: READ <= 8'Ha5;
		32'H00080001: READ <= 8'Ha7;
		32'H00080002: READ <= 8'Hab;
		32'H00080003: READ <= 8'Haf;
		32'H00080004: READ <= 8'Hb1;
		32'H00080005: READ <= 8'Hb5;
		32'H00080006: READ <= 8'Hb7;
		32'H00080007: READ <= 8'Hbb;
		32'H00080008: READ <= 8'Hbd;
		32'H00080009: READ <= 8'Hc1;
		32'H0008000a: READ <= 8'Hc5;
		32'H0008000b: READ <= 8'Hca;
		32'H0008000c: READ <= 8'Hcc;
		32'H0008000d: READ <= 8'Hd0;
		32'H0008000e: READ <= 8'Hd4;
		32'H0008000f: READ <= 8'Hd7;
		32'H00080010: READ <= 8'Hdb;
		32'H00080011: READ <= 8'Hde;
		32'H00080012: READ <= 8'He1;
		32'H00080013: READ <= 8'He4;
		32'H00080014: READ <= 8'He6;
		32'H00080015: READ <= 8'He9;
		32'H00080016: READ <= 8'Hea;
		32'H00080017: READ <= 8'Heb;
		32'H00080018: READ <= 8'Hed;
		32'H00080019: READ <= 8'Hee;
		32'H0008001a: READ <= 8'Hef;
		32'H0008001b: READ <= 8'Hf0;
		32'H0008001c: READ <= 8'Hf2;
		32'H0008001d: READ <= 8'Hf2;
		32'H0008001e: READ <= 8'Hf3;
		32'H0008001f: READ <= 8'Hf3;
		32'H00080020: READ <= 8'Hee;
		32'H00080021: READ <= 8'Hc2;
		32'H00080022: READ <= 8'H9c;
		32'H00080023: READ <= 8'H60;
		32'H00080024: READ <= 8'H62;
		32'H00080025: READ <= 8'H64;
		32'H00080026: READ <= 8'H7a;
		32'H00080027: READ <= 8'H83;
		32'H00080028: READ <= 8'H99;
		32'H00080029: READ <= 8'H97;
		32'H0008002a: READ <= 8'H98;
		32'H0008002b: READ <= 8'Haf;
		32'H0008002c: READ <= 8'H96;
		32'H0008002d: READ <= 8'H92;
		32'H0008002e: READ <= 8'H9a;
		32'H0008002f: READ <= 8'H9e;
		32'H00080030: READ <= 8'H81;
		32'H00080031: READ <= 8'H8b;
		32'H00080032: READ <= 8'H79;
		32'H00080033: READ <= 8'H8b;
		32'H00080034: READ <= 8'H82;
		32'H00080035: READ <= 8'H9a;
		32'H00080036: READ <= 8'H9e;
		32'H00080037: READ <= 8'Ha9;
		32'H00080038: READ <= 8'H9e;
		32'H00080039: READ <= 8'H99;
		32'H0008003a: READ <= 8'H98;
		32'H0008003b: READ <= 8'H96;
		32'H0008003c: READ <= 8'H95;
		32'H0008003d: READ <= 8'H93;
		32'H0008003e: READ <= 8'H91;
		32'H0008003f: READ <= 8'H91;
		32'H00080040: READ <= 8'H92;
		32'H00080041: READ <= 8'H92;
		32'H00080042: READ <= 8'H92;
		32'H00080043: READ <= 8'H93;
		32'H00080044: READ <= 8'H92;
		32'H00080045: READ <= 8'H93;
		32'H00080046: READ <= 8'H93;
		32'H00080047: READ <= 8'H94;
		32'H00080048: READ <= 8'H94;
		32'H00080049: READ <= 8'H95;
		32'H0008004a: READ <= 8'H94;
		32'H0008004b: READ <= 8'H96;
		32'H0008004c: READ <= 8'H95;
		32'H0008004d: READ <= 8'H96;
		32'H0008004e: READ <= 8'H98;
		32'H0008004f: READ <= 8'H99;
		32'H00080050: READ <= 8'H99;
		32'H00080051: READ <= 8'H99;
		32'H00080052: READ <= 8'H9a;
		32'H00080053: READ <= 8'H9b;
		32'H00080054: READ <= 8'H9b;
		32'H00080055: READ <= 8'H9c;
		32'H00080056: READ <= 8'H9d;
		32'H00080057: READ <= 8'H9c;
		32'H00080058: READ <= 8'H9c;
		32'H00080059: READ <= 8'H9c;
		32'H0008005a: READ <= 8'H9c;
		32'H0008005b: READ <= 8'H9d;
		32'H0008005c: READ <= 8'H9d;
		32'H0008005d: READ <= 8'H9c;
		32'H0008005e: READ <= 8'H9d;
		32'H0008005f: READ <= 8'H9c;
		32'H00080060: READ <= 8'H9d;
		32'H00080061: READ <= 8'H9e;
		32'H00080062: READ <= 8'H9e;
		32'H00080063: READ <= 8'H9f;
		
		32'H00090000: READ <= 8'Ha4;
		32'H00090001: READ <= 8'Ha7;
		32'H00090002: READ <= 8'Ha9;
		32'H00090003: READ <= 8'Had;
		32'H00090004: READ <= 8'Hb0;
		32'H00090005: READ <= 8'Hb3;
		32'H00090006: READ <= 8'Hb5;
		32'H00090007: READ <= 8'Hb9;
		32'H00090008: READ <= 8'Hbb;
		32'H00090009: READ <= 8'Hbf;
		32'H0009000a: READ <= 8'Hc3;
		32'H0009000b: READ <= 8'Hc7;
		32'H0009000c: READ <= 8'Hcb;
		32'H0009000d: READ <= 8'Hcf;
		32'H0009000e: READ <= 8'Hd2;
		32'H0009000f: READ <= 8'Hd6;
		32'H00090010: READ <= 8'Hd9;
		32'H00090011: READ <= 8'Hdd;
		32'H00090012: READ <= 8'He0;
		32'H00090013: READ <= 8'He4;
		32'H00090014: READ <= 8'He6;
		32'H00090015: READ <= 8'He7;
		32'H00090016: READ <= 8'Hea;
		32'H00090017: READ <= 8'Hec;
		32'H00090018: READ <= 8'Hed;
		32'H00090019: READ <= 8'Hed;
		32'H0009001a: READ <= 8'Hf0;
		32'H0009001b: READ <= 8'Hf1;
		32'H0009001c: READ <= 8'Hf1;
		32'H0009001d: READ <= 8'Hf3;
		32'H0009001e: READ <= 8'Hf1;
		32'H0009001f: READ <= 8'Hcb;
		32'H00090020: READ <= 8'Ha5;
		32'H00090021: READ <= 8'H88;
		32'H00090022: READ <= 8'H75;
		32'H00090023: READ <= 8'H81;
		32'H00090024: READ <= 8'H8c;
		32'H00090025: READ <= 8'H4a;
		32'H00090026: READ <= 8'H5f;
		32'H00090027: READ <= 8'Ha1;
		32'H00090028: READ <= 8'Ha6;
		32'H00090029: READ <= 8'H90;
		32'H0009002a: READ <= 8'H93;
		32'H0009002b: READ <= 8'H96;
		32'H0009002c: READ <= 8'H93;
		32'H0009002d: READ <= 8'H96;
		32'H0009002e: READ <= 8'H9e;
		32'H0009002f: READ <= 8'Hb1;
		32'H00090030: READ <= 8'H67;
		32'H00090031: READ <= 8'H7f;
		32'H00090032: READ <= 8'Hb0;
		32'H00090033: READ <= 8'Hc2;
		32'H00090034: READ <= 8'Hd8;
		32'H00090035: READ <= 8'Hdb;
		32'H00090036: READ <= 8'Hbd;
		32'H00090037: READ <= 8'Ha9;
		32'H00090038: READ <= 8'Hac;
		32'H00090039: READ <= 8'H9f;
		32'H0009003a: READ <= 8'H99;
		32'H0009003b: READ <= 8'H96;
		32'H0009003c: READ <= 8'H95;
		32'H0009003d: READ <= 8'H93;
		32'H0009003e: READ <= 8'H91;
		32'H0009003f: READ <= 8'H90;
		32'H00090040: READ <= 8'H90;
		32'H00090041: READ <= 8'H90;
		32'H00090042: READ <= 8'H91;
		32'H00090043: READ <= 8'H92;
		32'H00090044: READ <= 8'H92;
		32'H00090045: READ <= 8'H92;
		32'H00090046: READ <= 8'H92;
		32'H00090047: READ <= 8'H92;
		32'H00090048: READ <= 8'H92;
		32'H00090049: READ <= 8'H93;
		32'H0009004a: READ <= 8'H93;
		32'H0009004b: READ <= 8'H95;
		32'H0009004c: READ <= 8'H95;
		32'H0009004d: READ <= 8'H95;
		32'H0009004e: READ <= 8'H97;
		32'H0009004f: READ <= 8'H99;
		32'H00090050: READ <= 8'H98;
		32'H00090051: READ <= 8'H99;
		32'H00090052: READ <= 8'H9a;
		32'H00090053: READ <= 8'H9a;
		32'H00090054: READ <= 8'H9a;
		32'H00090055: READ <= 8'H9a;
		32'H00090056: READ <= 8'H9b;
		32'H00090057: READ <= 8'H9b;
		32'H00090058: READ <= 8'H9c;
		32'H00090059: READ <= 8'H9c;
		32'H0009005a: READ <= 8'H9b;
		32'H0009005b: READ <= 8'H9c;
		32'H0009005c: READ <= 8'H9b;
		32'H0009005d: READ <= 8'H9c;
		32'H0009005e: READ <= 8'H9c;
		32'H0009005f: READ <= 8'H9c;
		32'H00090060: READ <= 8'H9d;
		32'H00090061: READ <= 8'H9d;
		32'H00090062: READ <= 8'H9d;
		32'H00090063: READ <= 8'H9e;
		
		32'H000a0000: READ <= 8'Ha3;
		32'H000a0001: READ <= 8'Ha5;
		32'H000a0002: READ <= 8'Ha8;
		32'H000a0003: READ <= 8'Hab;
		32'H000a0004: READ <= 8'Hae;
		32'H000a0005: READ <= 8'Hb1;
		32'H000a0006: READ <= 8'Hb5;
		32'H000a0007: READ <= 8'Hb6;
		32'H000a0008: READ <= 8'Hba;
		32'H000a0009: READ <= 8'Hbd;
		32'H000a000a: READ <= 8'Hc0;
		32'H000a000b: READ <= 8'Hc5;
		32'H000a000c: READ <= 8'Hc9;
		32'H000a000d: READ <= 8'Hcd;
		32'H000a000e: READ <= 8'Hcf;
		32'H000a000f: READ <= 8'Hd3;
		32'H000a0010: READ <= 8'Hd7;
		32'H000a0011: READ <= 8'Hdb;
		32'H000a0012: READ <= 8'Hdf;
		32'H000a0013: READ <= 8'He2;
		32'H000a0014: READ <= 8'He4;
		32'H000a0015: READ <= 8'He7;
		32'H000a0016: READ <= 8'He9;
		32'H000a0017: READ <= 8'Heb;
		32'H000a0018: READ <= 8'Hec;
		32'H000a0019: READ <= 8'Hed;
		32'H000a001a: READ <= 8'Hef;
		32'H000a001b: READ <= 8'Hf2;
		32'H000a001c: READ <= 8'Hf2;
		32'H000a001d: READ <= 8'He6;
		32'H000a001e: READ <= 8'Haf;
		32'H000a001f: READ <= 8'H92;
		32'H000a0020: READ <= 8'H7f;
		32'H000a0021: READ <= 8'H8c;
		32'H000a0022: READ <= 8'H90;
		32'H000a0023: READ <= 8'H8a;
		32'H000a0024: READ <= 8'H8b;
		32'H000a0025: READ <= 8'H85;
		32'H000a0026: READ <= 8'H33;
		32'H000a0027: READ <= 8'H76;
		32'H000a0028: READ <= 8'H8e;
		32'H000a0029: READ <= 8'H96;
		32'H000a002a: READ <= 8'H81;
		32'H000a002b: READ <= 8'H88;
		32'H000a002c: READ <= 8'H97;
		32'H000a002d: READ <= 8'Ha3;
		32'H000a002e: READ <= 8'Hae;
		32'H000a002f: READ <= 8'H7a;
		32'H000a0030: READ <= 8'H9f;
		32'H000a0031: READ <= 8'Hc9;
		32'H000a0032: READ <= 8'Hd5;
		32'H000a0033: READ <= 8'Hde;
		32'H000a0034: READ <= 8'Hde;
		32'H000a0035: READ <= 8'Hda;
		32'H000a0036: READ <= 8'Hc1;
		32'H000a0037: READ <= 8'Haa;
		32'H000a0038: READ <= 8'Had;
		32'H000a0039: READ <= 8'H9a;
		32'H000a003a: READ <= 8'Ha0;
		32'H000a003b: READ <= 8'H9b;
		32'H000a003c: READ <= 8'H96;
		32'H000a003d: READ <= 8'H93;
		32'H000a003e: READ <= 8'H91;
		32'H000a003f: READ <= 8'H8f;
		32'H000a0040: READ <= 8'H8f;
		32'H000a0041: READ <= 8'H8e;
		32'H000a0042: READ <= 8'H90;
		32'H000a0043: READ <= 8'H90;
		32'H000a0044: READ <= 8'H91;
		32'H000a0045: READ <= 8'H91;
		32'H000a0046: READ <= 8'H90;
		32'H000a0047: READ <= 8'H92;
		32'H000a0048: READ <= 8'H92;
		32'H000a0049: READ <= 8'H91;
		32'H000a004a: READ <= 8'H93;
		32'H000a004b: READ <= 8'H93;
		32'H000a004c: READ <= 8'H94;
		32'H000a004d: READ <= 8'H96;
		32'H000a004e: READ <= 8'H97;
		32'H000a004f: READ <= 8'H97;
		32'H000a0050: READ <= 8'H98;
		32'H000a0051: READ <= 8'H98;
		32'H000a0052: READ <= 8'H98;
		32'H000a0053: READ <= 8'H99;
		32'H000a0054: READ <= 8'H99;
		32'H000a0055: READ <= 8'H99;
		32'H000a0056: READ <= 8'H99;
		32'H000a0057: READ <= 8'H9b;
		32'H000a0058: READ <= 8'H9b;
		32'H000a0059: READ <= 8'H9a;
		32'H000a005a: READ <= 8'H9a;
		32'H000a005b: READ <= 8'H9b;
		32'H000a005c: READ <= 8'H9b;
		32'H000a005d: READ <= 8'H9a;
		32'H000a005e: READ <= 8'H9a;
		32'H000a005f: READ <= 8'H9b;
		32'H000a0060: READ <= 8'H9b;
		32'H000a0061: READ <= 8'H9c;
		32'H000a0062: READ <= 8'H9c;
		32'H000a0063: READ <= 8'H9d;
		
		32'H000b0000: READ <= 8'Ha1;
		32'H000b0001: READ <= 8'Ha3;
		32'H000b0002: READ <= 8'Ha6;
		32'H000b0003: READ <= 8'Ha9;
		32'H000b0004: READ <= 8'Had;
		32'H000b0005: READ <= 8'Hb0;
		32'H000b0006: READ <= 8'Hb2;
		32'H000b0007: READ <= 8'Hb4;
		32'H000b0008: READ <= 8'Hb8;
		32'H000b0009: READ <= 8'Hbc;
		32'H000b000a: READ <= 8'Hbe;
		32'H000b000b: READ <= 8'Hc2;
		32'H000b000c: READ <= 8'Hc7;
		32'H000b000d: READ <= 8'Hcb;
		32'H000b000e: READ <= 8'Hcd;
		32'H000b000f: READ <= 8'Hd1;
		32'H000b0010: READ <= 8'Hd6;
		32'H000b0011: READ <= 8'Hd9;
		32'H000b0012: READ <= 8'Hdc;
		32'H000b0013: READ <= 8'He0;
		32'H000b0014: READ <= 8'He4;
		32'H000b0015: READ <= 8'He6;
		32'H000b0016: READ <= 8'He9;
		32'H000b0017: READ <= 8'Heb;
		32'H000b0018: READ <= 8'Hec;
		32'H000b0019: READ <= 8'Hed;
		32'H000b001a: READ <= 8'Hef;
		32'H000b001b: READ <= 8'Hf2;
		32'H000b001c: READ <= 8'Hd8;
		32'H000b001d: READ <= 8'Ha4;
		32'H000b001e: READ <= 8'H8e;
		32'H000b001f: READ <= 8'H87;
		32'H000b0020: READ <= 8'H91;
		32'H000b0021: READ <= 8'H9d;
		32'H000b0022: READ <= 8'H9c;
		32'H000b0023: READ <= 8'Ha0;
		32'H000b0024: READ <= 8'H98;
		32'H000b0025: READ <= 8'Ha6;
		32'H000b0026: READ <= 8'H81;
		32'H000b0027: READ <= 8'H88;
		32'H000b0028: READ <= 8'H97;
		32'H000b0029: READ <= 8'H76;
		32'H000b002a: READ <= 8'H65;
		32'H000b002b: READ <= 8'H82;
		32'H000b002c: READ <= 8'H9e;
		32'H000b002d: READ <= 8'Ha8;
		32'H000b002e: READ <= 8'Had;
		32'H000b002f: READ <= 8'Hc3;
		32'H000b0030: READ <= 8'Hcd;
		32'H000b0031: READ <= 8'Hd0;
		32'H000b0032: READ <= 8'Hd1;
		32'H000b0033: READ <= 8'Hcb;
		32'H000b0034: READ <= 8'Hc3;
		32'H000b0035: READ <= 8'Hba;
		32'H000b0036: READ <= 8'Hc2;
		32'H000b0037: READ <= 8'Hcc;
		32'H000b0038: READ <= 8'Hca;
		32'H000b0039: READ <= 8'Hac;
		32'H000b003a: READ <= 8'H96;
		32'H000b003b: READ <= 8'Ha5;
		32'H000b003c: READ <= 8'H9b;
		32'H000b003d: READ <= 8'H98;
		32'H000b003e: READ <= 8'H92;
		32'H000b003f: READ <= 8'H8e;
		32'H000b0040: READ <= 8'H8e;
		32'H000b0041: READ <= 8'H8e;
		32'H000b0042: READ <= 8'H8e;
		32'H000b0043: READ <= 8'H8f;
		32'H000b0044: READ <= 8'H8e;
		32'H000b0045: READ <= 8'H8f;
		32'H000b0046: READ <= 8'H8f;
		32'H000b0047: READ <= 8'H90;
		32'H000b0048: READ <= 8'H91;
		32'H000b0049: READ <= 8'H91;
		32'H000b004a: READ <= 8'H91;
		32'H000b004b: READ <= 8'H92;
		32'H000b004c: READ <= 8'H93;
		32'H000b004d: READ <= 8'H95;
		32'H000b004e: READ <= 8'H96;
		32'H000b004f: READ <= 8'H96;
		32'H000b0050: READ <= 8'H97;
		32'H000b0051: READ <= 8'H97;
		32'H000b0052: READ <= 8'H97;
		32'H000b0053: READ <= 8'H98;
		32'H000b0054: READ <= 8'H97;
		32'H000b0055: READ <= 8'H98;
		32'H000b0056: READ <= 8'H98;
		32'H000b0057: READ <= 8'H98;
		32'H000b0058: READ <= 8'H99;
		32'H000b0059: READ <= 8'H99;
		32'H000b005a: READ <= 8'H99;
		32'H000b005b: READ <= 8'H99;
		32'H000b005c: READ <= 8'H9a;
		32'H000b005d: READ <= 8'H9a;
		32'H000b005e: READ <= 8'H9a;
		32'H000b005f: READ <= 8'H99;
		32'H000b0060: READ <= 8'H99;
		32'H000b0061: READ <= 8'H9a;
		32'H000b0062: READ <= 8'H9a;
		32'H000b0063: READ <= 8'H9b;
		
		32'H000c0000: READ <= 8'H9f;
		32'H000c0001: READ <= 8'Ha2;
		32'H000c0002: READ <= 8'Ha4;
		32'H000c0003: READ <= 8'Ha7;
		32'H000c0004: READ <= 8'Hab;
		32'H000c0005: READ <= 8'Hae;
		32'H000c0006: READ <= 8'Hb1;
		32'H000c0007: READ <= 8'Hb3;
		32'H000c0008: READ <= 8'Hb7;
		32'H000c0009: READ <= 8'Hba;
		32'H000c000a: READ <= 8'Hbd;
		32'H000c000b: READ <= 8'Hc0;
		32'H000c000c: READ <= 8'Hc4;
		32'H000c000d: READ <= 8'Hc9;
		32'H000c000e: READ <= 8'Hcc;
		32'H000c000f: READ <= 8'Hce;
		32'H000c0010: READ <= 8'Hd2;
		32'H000c0011: READ <= 8'Hd6;
		32'H000c0012: READ <= 8'Hda;
		32'H000c0013: READ <= 8'Hdf;
		32'H000c0014: READ <= 8'He2;
		32'H000c0015: READ <= 8'He5;
		32'H000c0016: READ <= 8'He8;
		32'H000c0017: READ <= 8'Hea;
		32'H000c0018: READ <= 8'Hec;
		32'H000c0019: READ <= 8'Hee;
		32'H000c001a: READ <= 8'Hec;
		32'H000c001b: READ <= 8'Hd8;
		32'H000c001c: READ <= 8'Ha9;
		32'H000c001d: READ <= 8'H87;
		32'H000c001e: READ <= 8'H87;
		32'H000c001f: READ <= 8'H83;
		32'H000c0020: READ <= 8'H8c;
		32'H000c0021: READ <= 8'H9b;
		32'H000c0022: READ <= 8'H9a;
		32'H000c0023: READ <= 8'H9f;
		32'H000c0024: READ <= 8'Ha3;
		32'H000c0025: READ <= 8'H99;
		32'H000c0026: READ <= 8'Hab;
		32'H000c0027: READ <= 8'H9c;
		32'H000c0028: READ <= 8'H8b;
		32'H000c0029: READ <= 8'H5a;
		32'H000c002a: READ <= 8'H40;
		32'H000c002b: READ <= 8'H72;
		32'H000c002c: READ <= 8'Ha7;
		32'H000c002d: READ <= 8'Hb0;
		32'H000c002e: READ <= 8'Hc8;
		32'H000c002f: READ <= 8'Hd8;
		32'H000c0030: READ <= 8'Hd6;
		32'H000c0031: READ <= 8'Hc0;
		32'H000c0032: READ <= 8'Hb5;
		32'H000c0033: READ <= 8'Hb9;
		32'H000c0034: READ <= 8'Hc7;
		32'H000c0035: READ <= 8'Hd8;
		32'H000c0036: READ <= 8'Hd8;
		32'H000c0037: READ <= 8'Hda;
		32'H000c0038: READ <= 8'Hd3;
		32'H000c0039: READ <= 8'Hcf;
		32'H000c003a: READ <= 8'Hba;
		32'H000c003b: READ <= 8'H9c;
		32'H000c003c: READ <= 8'H9f;
		32'H000c003d: READ <= 8'H96;
		32'H000c003e: READ <= 8'H96;
		32'H000c003f: READ <= 8'H93;
		32'H000c0040: READ <= 8'H8d;
		32'H000c0041: READ <= 8'H8d;
		32'H000c0042: READ <= 8'H8d;
		32'H000c0043: READ <= 8'H8e;
		32'H000c0044: READ <= 8'H8d;
		32'H000c0045: READ <= 8'H8e;
		32'H000c0046: READ <= 8'H8f;
		32'H000c0047: READ <= 8'H8f;
		32'H000c0048: READ <= 8'H8f;
		32'H000c0049: READ <= 8'H90;
		32'H000c004a: READ <= 8'H91;
		32'H000c004b: READ <= 8'H91;
		32'H000c004c: READ <= 8'H92;
		32'H000c004d: READ <= 8'H93;
		32'H000c004e: READ <= 8'H96;
		32'H000c004f: READ <= 8'H96;
		32'H000c0050: READ <= 8'H96;
		32'H000c0051: READ <= 8'H96;
		32'H000c0052: READ <= 8'H97;
		32'H000c0053: READ <= 8'H97;
		32'H000c0054: READ <= 8'H97;
		32'H000c0055: READ <= 8'H97;
		32'H000c0056: READ <= 8'H97;
		32'H000c0057: READ <= 8'H97;
		32'H000c0058: READ <= 8'H97;
		32'H000c0059: READ <= 8'H97;
		32'H000c005a: READ <= 8'H98;
		32'H000c005b: READ <= 8'H98;
		32'H000c005c: READ <= 8'H99;
		32'H000c005d: READ <= 8'H99;
		32'H000c005e: READ <= 8'H99;
		32'H000c005f: READ <= 8'H98;
		32'H000c0060: READ <= 8'H99;
		32'H000c0061: READ <= 8'H99;
		32'H000c0062: READ <= 8'H99;
		32'H000c0063: READ <= 8'H9a;
		
		32'H000d0000: READ <= 8'H9e;
		32'H000d0001: READ <= 8'Ha0;
		32'H000d0002: READ <= 8'Ha2;
		32'H000d0003: READ <= 8'Ha5;
		32'H000d0004: READ <= 8'Haa;
		32'H000d0005: READ <= 8'Had;
		32'H000d0006: READ <= 8'Haf;
		32'H000d0007: READ <= 8'Hb2;
		32'H000d0008: READ <= 8'Hb5;
		32'H000d0009: READ <= 8'Hb8;
		32'H000d000a: READ <= 8'Hbb;
		32'H000d000b: READ <= 8'Hbe;
		32'H000d000c: READ <= 8'Hc1;
		32'H000d000d: READ <= 8'Hc6;
		32'H000d000e: READ <= 8'Hca;
		32'H000d000f: READ <= 8'Hcd;
		32'H000d0010: READ <= 8'Hcf;
		32'H000d0011: READ <= 8'Hd3;
		32'H000d0012: READ <= 8'Hd9;
		32'H000d0013: READ <= 8'Hdd;
		32'H000d0014: READ <= 8'He1;
		32'H000d0015: READ <= 8'He5;
		32'H000d0016: READ <= 8'He7;
		32'H000d0017: READ <= 8'He9;
		32'H000d0018: READ <= 8'Hec;
		32'H000d0019: READ <= 8'Hed;
		32'H000d001a: READ <= 8'Hd9;
		32'H000d001b: READ <= 8'Ha8;
		32'H000d001c: READ <= 8'H9e;
		32'H000d001d: READ <= 8'H8c;
		32'H000d001e: READ <= 8'H82;
		32'H000d001f: READ <= 8'H89;
		32'H000d0020: READ <= 8'H95;
		32'H000d0021: READ <= 8'H95;
		32'H000d0022: READ <= 8'H99;
		32'H000d0023: READ <= 8'H90;
		32'H000d0024: READ <= 8'H9c;
		32'H000d0025: READ <= 8'H93;
		32'H000d0026: READ <= 8'H92;
		32'H000d0027: READ <= 8'H73;
		32'H000d0028: READ <= 8'H5a;
		32'H000d0029: READ <= 8'H2d;
		32'H000d002a: READ <= 8'H20;
		32'H000d002b: READ <= 8'H67;
		32'H000d002c: READ <= 8'Ha4;
		32'H000d002d: READ <= 8'Hbd;
		32'H000d002e: READ <= 8'Hcf;
		32'H000d002f: READ <= 8'Hbd;
		32'H000d0030: READ <= 8'Hab;
		32'H000d0031: READ <= 8'Hb0;
		32'H000d0032: READ <= 8'Hc4;
		32'H000d0033: READ <= 8'Hd9;
		32'H000d0034: READ <= 8'Hd5;
		32'H000d0035: READ <= 8'Hdd;
		32'H000d0036: READ <= 8'Hdd;
		32'H000d0037: READ <= 8'Hd7;
		32'H000d0038: READ <= 8'Hce;
		32'H000d0039: READ <= 8'Hc1;
		32'H000d003a: READ <= 8'Hba;
		32'H000d003b: READ <= 8'Haf;
		32'H000d003c: READ <= 8'Ha5;
		32'H000d003d: READ <= 8'H97;
		32'H000d003e: READ <= 8'H8d;
		32'H000d003f: READ <= 8'H8e;
		32'H000d0040: READ <= 8'H95;
		32'H000d0041: READ <= 8'H93;
		32'H000d0042: READ <= 8'H8d;
		32'H000d0043: READ <= 8'H8c;
		32'H000d0044: READ <= 8'H8d;
		32'H000d0045: READ <= 8'H8c;
		32'H000d0046: READ <= 8'H8d;
		32'H000d0047: READ <= 8'H8e;
		32'H000d0048: READ <= 8'H8e;
		32'H000d0049: READ <= 8'H8f;
		32'H000d004a: READ <= 8'H90;
		32'H000d004b: READ <= 8'H91;
		32'H000d004c: READ <= 8'H91;
		32'H000d004d: READ <= 8'H93;
		32'H000d004e: READ <= 8'H94;
		32'H000d004f: READ <= 8'H94;
		32'H000d0050: READ <= 8'H95;
		32'H000d0051: READ <= 8'H96;
		32'H000d0052: READ <= 8'H96;
		32'H000d0053: READ <= 8'H96;
		32'H000d0054: READ <= 8'H95;
		32'H000d0055: READ <= 8'H96;
		32'H000d0056: READ <= 8'H96;
		32'H000d0057: READ <= 8'H96;
		32'H000d0058: READ <= 8'H96;
		32'H000d0059: READ <= 8'H97;
		32'H000d005a: READ <= 8'H97;
		32'H000d005b: READ <= 8'H98;
		32'H000d005c: READ <= 8'H97;
		32'H000d005d: READ <= 8'H97;
		32'H000d005e: READ <= 8'H97;
		32'H000d005f: READ <= 8'H97;
		32'H000d0060: READ <= 8'H98;
		32'H000d0061: READ <= 8'H98;
		32'H000d0062: READ <= 8'H99;
		32'H000d0063: READ <= 8'H99;
		
		32'H000e0000: READ <= 8'H9e;
		32'H000e0001: READ <= 8'H9e;
		32'H000e0002: READ <= 8'Ha1;
		32'H000e0003: READ <= 8'Ha4;
		32'H000e0004: READ <= 8'Ha7;
		32'H000e0005: READ <= 8'Hab;
		32'H000e0006: READ <= 8'Hae;
		32'H000e0007: READ <= 8'Hb0;
		32'H000e0008: READ <= 8'Hb2;
		32'H000e0009: READ <= 8'Hb6;
		32'H000e000a: READ <= 8'Hb9;
		32'H000e000b: READ <= 8'Hbc;
		32'H000e000c: READ <= 8'Hc0;
		32'H000e000d: READ <= 8'Hc4;
		32'H000e000e: READ <= 8'Hc8;
		32'H000e000f: READ <= 8'Hcb;
		32'H000e0010: READ <= 8'Hcd;
		32'H000e0011: READ <= 8'Hd0;
		32'H000e0012: READ <= 8'Hd5;
		32'H000e0013: READ <= 8'Hda;
		32'H000e0014: READ <= 8'He0;
		32'H000e0015: READ <= 8'He3;
		32'H000e0016: READ <= 8'He7;
		32'H000e0017: READ <= 8'He9;
		32'H000e0018: READ <= 8'Hec;
		32'H000e0019: READ <= 8'He8;
		32'H000e001a: READ <= 8'Hc0;
		32'H000e001b: READ <= 8'H99;
		32'H000e001c: READ <= 8'H95;
		32'H000e001d: READ <= 8'H82;
		32'H000e001e: READ <= 8'H92;
		32'H000e001f: READ <= 8'H93;
		32'H000e0020: READ <= 8'Ha0;
		32'H000e0021: READ <= 8'H97;
		32'H000e0022: READ <= 8'H94;
		32'H000e0023: READ <= 8'H94;
		32'H000e0024: READ <= 8'H8f;
		32'H000e0025: READ <= 8'H7f;
		32'H000e0026: READ <= 8'H70;
		32'H000e0027: READ <= 8'H2e;
		32'H000e0028: READ <= 8'H14;
		32'H000e0029: READ <= 8'H1a;
		32'H000e002a: READ <= 8'H41;
		32'H000e002b: READ <= 8'H8c;
		32'H000e002c: READ <= 8'H8f;
		32'H000e002d: READ <= 8'H97;
		32'H000e002e: READ <= 8'H97;
		32'H000e002f: READ <= 8'Ha2;
		32'H000e0030: READ <= 8'Hb8;
		32'H000e0031: READ <= 8'Hd0;
		32'H000e0032: READ <= 8'Hda;
		32'H000e0033: READ <= 8'He2;
		32'H000e0034: READ <= 8'Hd9;
		32'H000e0035: READ <= 8'Hc7;
		32'H000e0036: READ <= 8'Hbe;
		32'H000e0037: READ <= 8'Hc1;
		32'H000e0038: READ <= 8'Hca;
		32'H000e0039: READ <= 8'Hcc;
		32'H000e003a: READ <= 8'Hd1;
		32'H000e003b: READ <= 8'Hd4;
		32'H000e003c: READ <= 8'Hd0;
		32'H000e003d: READ <= 8'Hd0;
		32'H000e003e: READ <= 8'Had;
		32'H000e003f: READ <= 8'H9d;
		32'H000e0040: READ <= 8'H9b;
		32'H000e0041: READ <= 8'H93;
		32'H000e0042: READ <= 8'H95;
		32'H000e0043: READ <= 8'H8e;
		32'H000e0044: READ <= 8'H8a;
		32'H000e0045: READ <= 8'H8b;
		32'H000e0046: READ <= 8'H8b;
		32'H000e0047: READ <= 8'H8c;
		32'H000e0048: READ <= 8'H8d;
		32'H000e0049: READ <= 8'H8e;
		32'H000e004a: READ <= 8'H8f;
		32'H000e004b: READ <= 8'H8f;
		32'H000e004c: READ <= 8'H8f;
		32'H000e004d: READ <= 8'H91;
		32'H000e004e: READ <= 8'H92;
		32'H000e004f: READ <= 8'H92;
		32'H000e0050: READ <= 8'H94;
		32'H000e0051: READ <= 8'H94;
		32'H000e0052: READ <= 8'H94;
		32'H000e0053: READ <= 8'H94;
		32'H000e0054: READ <= 8'H95;
		32'H000e0055: READ <= 8'H96;
		32'H000e0056: READ <= 8'H95;
		32'H000e0057: READ <= 8'H95;
		32'H000e0058: READ <= 8'H96;
		32'H000e0059: READ <= 8'H96;
		32'H000e005a: READ <= 8'H96;
		32'H000e005b: READ <= 8'H96;
		32'H000e005c: READ <= 8'H96;
		32'H000e005d: READ <= 8'H97;
		32'H000e005e: READ <= 8'H97;
		32'H000e005f: READ <= 8'H96;
		32'H000e0060: READ <= 8'H97;
		32'H000e0061: READ <= 8'H97;
		32'H000e0062: READ <= 8'H97;
		32'H000e0063: READ <= 8'H97;
		
		32'H000f0000: READ <= 8'H9c;
		32'H000f0001: READ <= 8'H9d;
		32'H000f0002: READ <= 8'Ha0;
		32'H000f0003: READ <= 8'Ha3;
		32'H000f0004: READ <= 8'Ha5;
		32'H000f0005: READ <= 8'Ha9;
		32'H000f0006: READ <= 8'Hac;
		32'H000f0007: READ <= 8'Haf;
		32'H000f0008: READ <= 8'Hb1;
		32'H000f0009: READ <= 8'Hb4;
		32'H000f000a: READ <= 8'Hb8;
		32'H000f000b: READ <= 8'Hbb;
		32'H000f000c: READ <= 8'Hbe;
		32'H000f000d: READ <= 8'Hc2;
		32'H000f000e: READ <= 8'Hc5;
		32'H000f000f: READ <= 8'Hc9;
		32'H000f0010: READ <= 8'Hcb;
		32'H000f0011: READ <= 8'Hcf;
		32'H000f0012: READ <= 8'Hd3;
		32'H000f0013: READ <= 8'Hd8;
		32'H000f0014: READ <= 8'Hdd;
		32'H000f0015: READ <= 8'He1;
		32'H000f0016: READ <= 8'He5;
		32'H000f0017: READ <= 8'Hea;
		32'H000f0018: READ <= 8'He9;
		32'H000f0019: READ <= 8'Hd2;
		32'H000f001a: READ <= 8'Haf;
		32'H000f001b: READ <= 8'Hab;
		32'H000f001c: READ <= 8'H98;
		32'H000f001d: READ <= 8'H89;
		32'H000f001e: READ <= 8'H92;
		32'H000f001f: READ <= 8'H90;
		32'H000f0020: READ <= 8'H98;
		32'H000f0021: READ <= 8'H89;
		32'H000f0022: READ <= 8'H7d;
		32'H000f0023: READ <= 8'H72;
		32'H000f0024: READ <= 8'H8a;
		32'H000f0025: READ <= 8'H62;
		32'H000f0026: READ <= 8'H34;
		32'H000f0027: READ <= 8'H1;
		32'H000f0028: READ <= 8'H16;
		32'H000f0029: READ <= 8'H5f;
		32'H000f002a: READ <= 8'H91;
		32'H000f002b: READ <= 8'Ha8;
		32'H000f002c: READ <= 8'H8f;
		32'H000f002d: READ <= 8'H82;
		32'H000f002e: READ <= 8'H9f;
		32'H000f002f: READ <= 8'Hcb;
		32'H000f0030: READ <= 8'Hcd;
		32'H000f0031: READ <= 8'Hc8;
		32'H000f0032: READ <= 8'Hbe;
		32'H000f0033: READ <= 8'Haf;
		32'H000f0034: READ <= 8'Had;
		32'H000f0035: READ <= 8'Hb3;
		32'H000f0036: READ <= 8'Hcf;
		32'H000f0037: READ <= 8'Hd9;
		32'H000f0038: READ <= 8'Hdc;
		32'H000f0039: READ <= 8'Hdf;
		32'H000f003a: READ <= 8'He8;
		32'H000f003b: READ <= 8'He7;
		32'H000f003c: READ <= 8'He0;
		32'H000f003d: READ <= 8'Hdd;
		32'H000f003e: READ <= 8'Hd7;
		32'H000f003f: READ <= 8'H9e;
		32'H000f0040: READ <= 8'H9a;
		32'H000f0041: READ <= 8'H91;
		32'H000f0042: READ <= 8'H87;
		32'H000f0043: READ <= 8'H8a;
		32'H000f0044: READ <= 8'H92;
		32'H000f0045: READ <= 8'H89;
		32'H000f0046: READ <= 8'H8a;
		32'H000f0047: READ <= 8'H8b;
		32'H000f0048: READ <= 8'H8c;
		32'H000f0049: READ <= 8'H8c;
		32'H000f004a: READ <= 8'H8e;
		32'H000f004b: READ <= 8'H8e;
		32'H000f004c: READ <= 8'H8f;
		32'H000f004d: READ <= 8'H8f;
		32'H000f004e: READ <= 8'H91;
		32'H000f004f: READ <= 8'H91;
		32'H000f0050: READ <= 8'H92;
		32'H000f0051: READ <= 8'H93;
		32'H000f0052: READ <= 8'H93;
		32'H000f0053: READ <= 8'H93;
		32'H000f0054: READ <= 8'H94;
		32'H000f0055: READ <= 8'H94;
		32'H000f0056: READ <= 8'H94;
		32'H000f0057: READ <= 8'H94;
		32'H000f0058: READ <= 8'H94;
		32'H000f0059: READ <= 8'H94;
		32'H000f005a: READ <= 8'H94;
		32'H000f005b: READ <= 8'H95;
		32'H000f005c: READ <= 8'H96;
		32'H000f005d: READ <= 8'H96;
		32'H000f005e: READ <= 8'H96;
		32'H000f005f: READ <= 8'H96;
		32'H000f0060: READ <= 8'H96;
		32'H000f0061: READ <= 8'H96;
		32'H000f0062: READ <= 8'H96;
		32'H000f0063: READ <= 8'H96;
		
		32'H00100000: READ <= 8'H9a;
		32'H00100001: READ <= 8'H9c;
		32'H00100002: READ <= 8'H9e;
		32'H00100003: READ <= 8'Ha0;
		32'H00100004: READ <= 8'Ha4;
		32'H00100005: READ <= 8'Ha7;
		32'H00100006: READ <= 8'Haa;
		32'H00100007: READ <= 8'Had;
		32'H00100008: READ <= 8'Hb0;
		32'H00100009: READ <= 8'Hb2;
		32'H0010000a: READ <= 8'Hb7;
		32'H0010000b: READ <= 8'Hba;
		32'H0010000c: READ <= 8'Hbc;
		32'H0010000d: READ <= 8'Hbe;
		32'H0010000e: READ <= 8'Hc3;
		32'H0010000f: READ <= 8'Hc7;
		32'H00100010: READ <= 8'Hc9;
		32'H00100011: READ <= 8'Hcd;
		32'H00100012: READ <= 8'Hd0;
		32'H00100013: READ <= 8'Hd6;
		32'H00100014: READ <= 8'Hdb;
		32'H00100015: READ <= 8'He0;
		32'H00100016: READ <= 8'He3;
		32'H00100017: READ <= 8'He6;
		32'H00100018: READ <= 8'He9;
		32'H00100019: READ <= 8'Hc7;
		32'H0010001a: READ <= 8'Haf;
		32'H0010001b: READ <= 8'Hb1;
		32'H0010001c: READ <= 8'H91;
		32'H0010001d: READ <= 8'H8d;
		32'H0010001e: READ <= 8'H9d;
		32'H0010001f: READ <= 8'H97;
		32'H00100020: READ <= 8'H96;
		32'H00100021: READ <= 8'H6d;
		32'H00100022: READ <= 8'H82;
		32'H00100023: READ <= 8'H6f;
		32'H00100024: READ <= 8'H70;
		32'H00100025: READ <= 8'H41;
		32'H00100026: READ <= 8'H0;
		32'H00100027: READ <= 8'H38;
		32'H00100028: READ <= 8'H8c;
		32'H00100029: READ <= 8'H97;
		32'H0010002a: READ <= 8'Ha8;
		32'H0010002b: READ <= 8'H88;
		32'H0010002c: READ <= 8'H86;
		32'H0010002d: READ <= 8'Hb3;
		32'H0010002e: READ <= 8'Hbd;
		32'H0010002f: READ <= 8'Hc3;
		32'H00100030: READ <= 8'Hb0;
		32'H00100031: READ <= 8'Had;
		32'H00100032: READ <= 8'Haa;
		32'H00100033: READ <= 8'Hb7;
		32'H00100034: READ <= 8'Hc8;
		32'H00100035: READ <= 8'Hd2;
		32'H00100036: READ <= 8'Hd8;
		32'H00100037: READ <= 8'Hd8;
		32'H00100038: READ <= 8'Hdc;
		32'H00100039: READ <= 8'He1;
		32'H0010003a: READ <= 8'He8;
		32'H0010003b: READ <= 8'Heb;
		32'H0010003c: READ <= 8'He7;
		32'H0010003d: READ <= 8'Hd9;
		32'H0010003e: READ <= 8'Hd5;
		32'H0010003f: READ <= 8'Hc2;
		32'H00100040: READ <= 8'H86;
		32'H00100041: READ <= 8'H82;
		32'H00100042: READ <= 8'H82;
		32'H00100043: READ <= 8'H7d;
		32'H00100044: READ <= 8'H88;
		32'H00100045: READ <= 8'H96;
		32'H00100046: READ <= 8'H8c;
		32'H00100047: READ <= 8'H8a;
		32'H00100048: READ <= 8'H8a;
		32'H00100049: READ <= 8'H8b;
		32'H0010004a: READ <= 8'H8c;
		32'H0010004b: READ <= 8'H8d;
		32'H0010004c: READ <= 8'H8d;
		32'H0010004d: READ <= 8'H8f;
		32'H0010004e: READ <= 8'H8f;
		32'H0010004f: READ <= 8'H90;
		32'H00100050: READ <= 8'H91;
		32'H00100051: READ <= 8'H92;
		32'H00100052: READ <= 8'H92;
		32'H00100053: READ <= 8'H92;
		32'H00100054: READ <= 8'H93;
		32'H00100055: READ <= 8'H92;
		32'H00100056: READ <= 8'H92;
		32'H00100057: READ <= 8'H93;
		32'H00100058: READ <= 8'H93;
		32'H00100059: READ <= 8'H93;
		32'H0010005a: READ <= 8'H94;
		32'H0010005b: READ <= 8'H94;
		32'H0010005c: READ <= 8'H94;
		32'H0010005d: READ <= 8'H95;
		32'H0010005e: READ <= 8'H95;
		32'H0010005f: READ <= 8'H95;
		32'H00100060: READ <= 8'H95;
		32'H00100061: READ <= 8'H95;
		32'H00100062: READ <= 8'H95;
		32'H00100063: READ <= 8'H95;
		
		32'H00110000: READ <= 8'H97;
		32'H00110001: READ <= 8'H9a;
		32'H00110002: READ <= 8'H9b;
		32'H00110003: READ <= 8'H9e;
		32'H00110004: READ <= 8'Ha1;
		32'H00110005: READ <= 8'Ha5;
		32'H00110006: READ <= 8'Ha8;
		32'H00110007: READ <= 8'Hab;
		32'H00110008: READ <= 8'Hae;
		32'H00110009: READ <= 8'Hb1;
		32'H0011000a: READ <= 8'Hb4;
		32'H0011000b: READ <= 8'Hb8;
		32'H0011000c: READ <= 8'Hbb;
		32'H0011000d: READ <= 8'Hbc;
		32'H0011000e: READ <= 8'Hc1;
		32'H0011000f: READ <= 8'Hc5;
		32'H00110010: READ <= 8'Hc7;
		32'H00110011: READ <= 8'Hca;
		32'H00110012: READ <= 8'Hcf;
		32'H00110013: READ <= 8'Hd4;
		32'H00110014: READ <= 8'Hd8;
		32'H00110015: READ <= 8'Hdd;
		32'H00110016: READ <= 8'He1;
		32'H00110017: READ <= 8'He4;
		32'H00110018: READ <= 8'He2;
		32'H00110019: READ <= 8'Hb1;
		32'H0011001a: READ <= 8'Hab;
		32'H0011001b: READ <= 8'Ha0;
		32'H0011001c: READ <= 8'H88;
		32'H0011001d: READ <= 8'H8f;
		32'H0011001e: READ <= 8'H9a;
		32'H0011001f: READ <= 8'H84;
		32'H00110020: READ <= 8'H77;
		32'H00110021: READ <= 8'H7a;
		32'H00110022: READ <= 8'H71;
		32'H00110023: READ <= 8'H73;
		32'H00110024: READ <= 8'H57;
		32'H00110025: READ <= 8'H26;
		32'H00110026: READ <= 8'H2a;
		32'H00110027: READ <= 8'H7e;
		32'H00110028: READ <= 8'H79;
		32'H00110029: READ <= 8'H8e;
		32'H0011002a: READ <= 8'Ha2;
		32'H0011002b: READ <= 8'H7f;
		32'H0011002c: READ <= 8'H63;
		32'H0011002d: READ <= 8'H80;
		32'H0011002e: READ <= 8'H9d;
		32'H0011002f: READ <= 8'H7c;
		32'H00110030: READ <= 8'H85;
		32'H00110031: READ <= 8'H91;
		32'H00110032: READ <= 8'Ha3;
		32'H00110033: READ <= 8'Ha4;
		32'H00110034: READ <= 8'Haa;
		32'H00110035: READ <= 8'Hb0;
		32'H00110036: READ <= 8'Hb6;
		32'H00110037: READ <= 8'Hb4;
		32'H00110038: READ <= 8'Hb8;
		32'H00110039: READ <= 8'Hc0;
		32'H0011003a: READ <= 8'Hc6;
		32'H0011003b: READ <= 8'Hce;
		32'H0011003c: READ <= 8'Hc7;
		32'H0011003d: READ <= 8'Hbc;
		32'H0011003e: READ <= 8'Hbe;
		32'H0011003f: READ <= 8'Hcd;
		32'H00110040: READ <= 8'Hc5;
		32'H00110041: READ <= 8'H9c;
		32'H00110042: READ <= 8'H7f;
		32'H00110043: READ <= 8'H8c;
		32'H00110044: READ <= 8'H75;
		32'H00110045: READ <= 8'H83;
		32'H00110046: READ <= 8'H93;
		32'H00110047: READ <= 8'H8e;
		32'H00110048: READ <= 8'H88;
		32'H00110049: READ <= 8'H89;
		32'H0011004a: READ <= 8'H8b;
		32'H0011004b: READ <= 8'H8b;
		32'H0011004c: READ <= 8'H8c;
		32'H0011004d: READ <= 8'H8d;
		32'H0011004e: READ <= 8'H8e;
		32'H0011004f: READ <= 8'H8f;
		32'H00110050: READ <= 8'H8f;
		32'H00110051: READ <= 8'H90;
		32'H00110052: READ <= 8'H92;
		32'H00110053: READ <= 8'H92;
		32'H00110054: READ <= 8'H92;
		32'H00110055: READ <= 8'H91;
		32'H00110056: READ <= 8'H91;
		32'H00110057: READ <= 8'H92;
		32'H00110058: READ <= 8'H93;
		32'H00110059: READ <= 8'H93;
		32'H0011005a: READ <= 8'H93;
		32'H0011005b: READ <= 8'H94;
		32'H0011005c: READ <= 8'H93;
		32'H0011005d: READ <= 8'H94;
		32'H0011005e: READ <= 8'H94;
		32'H0011005f: READ <= 8'H94;
		32'H00110060: READ <= 8'H95;
		32'H00110061: READ <= 8'H94;
		32'H00110062: READ <= 8'H94;
		32'H00110063: READ <= 8'H95;
		
		32'H00120000: READ <= 8'H95;
		32'H00120001: READ <= 8'H97;
		32'H00120002: READ <= 8'H99;
		32'H00120003: READ <= 8'H9b;
		32'H00120004: READ <= 8'H9f;
		32'H00120005: READ <= 8'Ha3;
		32'H00120006: READ <= 8'Ha6;
		32'H00120007: READ <= 8'Ha9;
		32'H00120008: READ <= 8'Hac;
		32'H00120009: READ <= 8'Haf;
		32'H0012000a: READ <= 8'Hb3;
		32'H0012000b: READ <= 8'Hb6;
		32'H0012000c: READ <= 8'Hb9;
		32'H0012000d: READ <= 8'Hbb;
		32'H0012000e: READ <= 8'Hbf;
		32'H0012000f: READ <= 8'Hc3;
		32'H00120010: READ <= 8'Hc5;
		32'H00120011: READ <= 8'Hc8;
		32'H00120012: READ <= 8'Hcc;
		32'H00120013: READ <= 8'Hd0;
		32'H00120014: READ <= 8'Hd5;
		32'H00120015: READ <= 8'Hdb;
		32'H00120016: READ <= 8'Hde;
		32'H00120017: READ <= 8'He1;
		32'H00120018: READ <= 8'Hca;
		32'H00120019: READ <= 8'Ha9;
		32'H0012001a: READ <= 8'Ha3;
		32'H0012001b: READ <= 8'H9e;
		32'H0012001c: READ <= 8'H7c;
		32'H0012001d: READ <= 8'H7e;
		32'H0012001e: READ <= 8'H7b;
		32'H0012001f: READ <= 8'H87;
		32'H00120020: READ <= 8'H6c;
		32'H00120021: READ <= 8'H82;
		32'H00120022: READ <= 8'H82;
		32'H00120023: READ <= 8'H74;
		32'H00120024: READ <= 8'H5b;
		32'H00120025: READ <= 8'Ha;
		32'H00120026: READ <= 8'H4e;
		32'H00120027: READ <= 8'H50;
		32'H00120028: READ <= 8'H43;
		32'H00120029: READ <= 8'H4d;
		32'H0012002a: READ <= 8'H71;
		32'H0012002b: READ <= 8'H63;
		32'H0012002c: READ <= 8'H6d;
		32'H0012002d: READ <= 8'H3d;
		32'H0012002e: READ <= 8'H5e;
		32'H0012002f: READ <= 8'H76;
		32'H00120030: READ <= 8'H72;
		32'H00120031: READ <= 8'H70;
		32'H00120032: READ <= 8'H6c;
		32'H00120033: READ <= 8'H6e;
		32'H00120034: READ <= 8'H69;
		32'H00120035: READ <= 8'H62;
		32'H00120036: READ <= 8'H61;
		32'H00120037: READ <= 8'H64;
		32'H00120038: READ <= 8'H69;
		32'H00120039: READ <= 8'H6e;
		32'H0012003a: READ <= 8'H7a;
		32'H0012003b: READ <= 8'H90;
		32'H0012003c: READ <= 8'H90;
		32'H0012003d: READ <= 8'H95;
		32'H0012003e: READ <= 8'H95;
		32'H0012003f: READ <= 8'H93;
		32'H00120040: READ <= 8'H99;
		32'H00120041: READ <= 8'H9c;
		32'H00120042: READ <= 8'H9c;
		32'H00120043: READ <= 8'H94;
		32'H00120044: READ <= 8'H76;
		32'H00120045: READ <= 8'H72;
		32'H00120046: READ <= 8'H7b;
		32'H00120047: READ <= 8'H8e;
		32'H00120048: READ <= 8'H93;
		32'H00120049: READ <= 8'H8a;
		32'H0012004a: READ <= 8'H8a;
		32'H0012004b: READ <= 8'H8a;
		32'H0012004c: READ <= 8'H8c;
		32'H0012004d: READ <= 8'H8c;
		32'H0012004e: READ <= 8'H8d;
		32'H0012004f: READ <= 8'H8e;
		32'H00120050: READ <= 8'H8e;
		32'H00120051: READ <= 8'H8f;
		32'H00120052: READ <= 8'H8f;
		32'H00120053: READ <= 8'H90;
		32'H00120054: READ <= 8'H91;
		32'H00120055: READ <= 8'H90;
		32'H00120056: READ <= 8'H90;
		32'H00120057: READ <= 8'H90;
		32'H00120058: READ <= 8'H92;
		32'H00120059: READ <= 8'H93;
		32'H0012005a: READ <= 8'H92;
		32'H0012005b: READ <= 8'H93;
		32'H0012005c: READ <= 8'H93;
		32'H0012005d: READ <= 8'H93;
		32'H0012005e: READ <= 8'H93;
		32'H0012005f: READ <= 8'H94;
		32'H00120060: READ <= 8'H94;
		32'H00120061: READ <= 8'H93;
		32'H00120062: READ <= 8'H94;
		32'H00120063: READ <= 8'H94;
		
		32'H00130000: READ <= 8'H93;
		32'H00130001: READ <= 8'H94;
		32'H00130002: READ <= 8'H97;
		32'H00130003: READ <= 8'H99;
		32'H00130004: READ <= 8'H9c;
		32'H00130005: READ <= 8'Ha0;
		32'H00130006: READ <= 8'Ha4;
		32'H00130007: READ <= 8'Ha7;
		32'H00130008: READ <= 8'Haa;
		32'H00130009: READ <= 8'Hae;
		32'H0013000a: READ <= 8'Hb1;
		32'H0013000b: READ <= 8'Hb3;
		32'H0013000c: READ <= 8'Hb7;
		32'H0013000d: READ <= 8'Hbb;
		32'H0013000e: READ <= 8'Hbe;
		32'H0013000f: READ <= 8'Hc1;
		32'H00130010: READ <= 8'Hc4;
		32'H00130011: READ <= 8'Hc6;
		32'H00130012: READ <= 8'Hca;
		32'H00130013: READ <= 8'Hcd;
		32'H00130014: READ <= 8'Hd2;
		32'H00130015: READ <= 8'Hd7;
		32'H00130016: READ <= 8'Hdd;
		32'H00130017: READ <= 8'Hdd;
		32'H00130018: READ <= 8'Hb4;
		32'H00130019: READ <= 8'Ha7;
		32'H0013001a: READ <= 8'H9f;
		32'H0013001b: READ <= 8'H93;
		32'H0013001c: READ <= 8'H6c;
		32'H0013001d: READ <= 8'H7f;
		32'H0013001e: READ <= 8'H77;
		32'H0013001f: READ <= 8'H70;
		32'H00130020: READ <= 8'H7d;
		32'H00130021: READ <= 8'H7f;
		32'H00130022: READ <= 8'H6d;
		32'H00130023: READ <= 8'H76;
		32'H00130024: READ <= 8'H40;
		32'H00130025: READ <= 8'H17;
		32'H00130026: READ <= 8'H4c;
		32'H00130027: READ <= 8'H48;
		32'H00130028: READ <= 8'H2f;
		32'H00130029: READ <= 8'H31;
		32'H0013002a: READ <= 8'H3c;
		32'H0013002b: READ <= 8'H20;
		32'H0013002c: READ <= 8'H2c;
		32'H0013002d: READ <= 8'H44;
		32'H0013002e: READ <= 8'H4a;
		32'H0013002f: READ <= 8'H5e;
		32'H00130030: READ <= 8'H63;
		32'H00130031: READ <= 8'H5f;
		32'H00130032: READ <= 8'H59;
		32'H00130033: READ <= 8'H54;
		32'H00130034: READ <= 8'H51;
		32'H00130035: READ <= 8'H50;
		32'H00130036: READ <= 8'H58;
		32'H00130037: READ <= 8'H61;
		32'H00130038: READ <= 8'H6f;
		32'H00130039: READ <= 8'H81;
		32'H0013003a: READ <= 8'H8f;
		32'H0013003b: READ <= 8'H9b;
		32'H0013003c: READ <= 8'H98;
		32'H0013003d: READ <= 8'H96;
		32'H0013003e: READ <= 8'H96;
		32'H0013003f: READ <= 8'H9e;
		32'H00130040: READ <= 8'H9d;
		32'H00130041: READ <= 8'H8b;
		32'H00130042: READ <= 8'H74;
		32'H00130043: READ <= 8'H71;
		32'H00130044: READ <= 8'H76;
		32'H00130045: READ <= 8'H7f;
		32'H00130046: READ <= 8'H80;
		32'H00130047: READ <= 8'H7b;
		32'H00130048: READ <= 8'H8a;
		32'H00130049: READ <= 8'H97;
		32'H0013004a: READ <= 8'H8e;
		32'H0013004b: READ <= 8'H89;
		32'H0013004c: READ <= 8'H8a;
		32'H0013004d: READ <= 8'H8b;
		32'H0013004e: READ <= 8'H8c;
		32'H0013004f: READ <= 8'H8c;
		32'H00130050: READ <= 8'H8d;
		32'H00130051: READ <= 8'H8e;
		32'H00130052: READ <= 8'H8f;
		32'H00130053: READ <= 8'H8f;
		32'H00130054: READ <= 8'H8f;
		32'H00130055: READ <= 8'H8f;
		32'H00130056: READ <= 8'H8f;
		32'H00130057: READ <= 8'H90;
		32'H00130058: READ <= 8'H91;
		32'H00130059: READ <= 8'H91;
		32'H0013005a: READ <= 8'H92;
		32'H0013005b: READ <= 8'H92;
		32'H0013005c: READ <= 8'H92;
		32'H0013005d: READ <= 8'H92;
		32'H0013005e: READ <= 8'H93;
		32'H0013005f: READ <= 8'H93;
		32'H00130060: READ <= 8'H93;
		32'H00130061: READ <= 8'H93;
		32'H00130062: READ <= 8'H93;
		32'H00130063: READ <= 8'H93;
		
		32'H00140000: READ <= 8'H91;
		32'H00140001: READ <= 8'H93;
		32'H00140002: READ <= 8'H95;
		32'H00140003: READ <= 8'H97;
		32'H00140004: READ <= 8'H9a;
		32'H00140005: READ <= 8'H9d;
		32'H00140006: READ <= 8'Ha1;
		32'H00140007: READ <= 8'Ha5;
		32'H00140008: READ <= 8'Haa;
		32'H00140009: READ <= 8'Hac;
		32'H0014000a: READ <= 8'Haf;
		32'H0014000b: READ <= 8'Hb1;
		32'H0014000c: READ <= 8'Hb5;
		32'H0014000d: READ <= 8'Hba;
		32'H0014000e: READ <= 8'Hbc;
		32'H0014000f: READ <= 8'Hbf;
		32'H00140010: READ <= 8'Hc2;
		32'H00140011: READ <= 8'Hc4;
		32'H00140012: READ <= 8'Hc8;
		32'H00140013: READ <= 8'Hcb;
		32'H00140014: READ <= 8'Hd0;
		32'H00140015: READ <= 8'Hd5;
		32'H00140016: READ <= 8'Hda;
		32'H00140017: READ <= 8'Hcc;
		32'H00140018: READ <= 8'Hb3;
		32'H00140019: READ <= 8'Ha9;
		32'H0014001a: READ <= 8'H94;
		32'H0014001b: READ <= 8'H87;
		32'H0014001c: READ <= 8'H5d;
		32'H0014001d: READ <= 8'H7e;
		32'H0014001e: READ <= 8'H6e;
		32'H0014001f: READ <= 8'H70;
		32'H00140020: READ <= 8'H72;
		32'H00140021: READ <= 8'H71;
		32'H00140022: READ <= 8'H84;
		32'H00140023: READ <= 8'H7a;
		32'H00140024: READ <= 8'H42;
		32'H00140025: READ <= 8'H14;
		32'H00140026: READ <= 8'H42;
		32'H00140027: READ <= 8'H2c;
		32'H00140028: READ <= 8'H23;
		32'H00140029: READ <= 8'H31;
		32'H0014002a: READ <= 8'H25;
		32'H0014002b: READ <= 8'H19;
		32'H0014002c: READ <= 8'H24;
		32'H0014002d: READ <= 8'H21;
		32'H0014002e: READ <= 8'H1c;
		32'H0014002f: READ <= 8'H38;
		32'H00140030: READ <= 8'H43;
		32'H00140031: READ <= 8'H32;
		32'H00140032: READ <= 8'H2b;
		32'H00140033: READ <= 8'H31;
		32'H00140034: READ <= 8'H41;
		32'H00140035: READ <= 8'H3a;
		32'H00140036: READ <= 8'H2f;
		32'H00140037: READ <= 8'H36;
		32'H00140038: READ <= 8'H3a;
		32'H00140039: READ <= 8'H3f;
		32'H0014003a: READ <= 8'H48;
		32'H0014003b: READ <= 8'H48;
		32'H0014003c: READ <= 8'H54;
		32'H0014003d: READ <= 8'H4a;
		32'H0014003e: READ <= 8'H40;
		32'H0014003f: READ <= 8'H49;
		32'H00140040: READ <= 8'H53;
		32'H00140041: READ <= 8'H56;
		32'H00140042: READ <= 8'H44;
		32'H00140043: READ <= 8'H41;
		32'H00140044: READ <= 8'H47;
		32'H00140045: READ <= 8'H52;
		32'H00140046: READ <= 8'H64;
		32'H00140047: READ <= 8'H74;
		32'H00140048: READ <= 8'H79;
		32'H00140049: READ <= 8'H84;
		32'H0014004a: READ <= 8'H93;
		32'H0014004b: READ <= 8'H8e;
		32'H0014004c: READ <= 8'H89;
		32'H0014004d: READ <= 8'H89;
		32'H0014004e: READ <= 8'H8a;
		32'H0014004f: READ <= 8'H8b;
		32'H00140050: READ <= 8'H8c;
		32'H00140051: READ <= 8'H8d;
		32'H00140052: READ <= 8'H8d;
		32'H00140053: READ <= 8'H8e;
		32'H00140054: READ <= 8'H8d;
		32'H00140055: READ <= 8'H8d;
		32'H00140056: READ <= 8'H8d;
		32'H00140057: READ <= 8'H8e;
		32'H00140058: READ <= 8'H8f;
		32'H00140059: READ <= 8'H90;
		32'H0014005a: READ <= 8'H90;
		32'H0014005b: READ <= 8'H91;
		32'H0014005c: READ <= 8'H92;
		32'H0014005d: READ <= 8'H92;
		32'H0014005e: READ <= 8'H92;
		32'H0014005f: READ <= 8'H92;
		32'H00140060: READ <= 8'H91;
		32'H00140061: READ <= 8'H92;
		32'H00140062: READ <= 8'H91;
		32'H00140063: READ <= 8'H91;
		
		32'H00150000: READ <= 8'H90;
		32'H00150001: READ <= 8'H91;
		32'H00150002: READ <= 8'H93;
		32'H00150003: READ <= 8'H95;
		32'H00150004: READ <= 8'H97;
		32'H00150005: READ <= 8'H9a;
		32'H00150006: READ <= 8'H9e;
		32'H00150007: READ <= 8'Ha2;
		32'H00150008: READ <= 8'Ha7;
		32'H00150009: READ <= 8'Hab;
		32'H0015000a: READ <= 8'Had;
		32'H0015000b: READ <= 8'Hb0;
		32'H0015000c: READ <= 8'Hb4;
		32'H0015000d: READ <= 8'Hb7;
		32'H0015000e: READ <= 8'Hbb;
		32'H0015000f: READ <= 8'Hbd;
		32'H00150010: READ <= 8'Hbf;
		32'H00150011: READ <= 8'Hc2;
		32'H00150012: READ <= 8'Hc5;
		32'H00150013: READ <= 8'Hc8;
		32'H00150014: READ <= 8'Hcd;
		32'H00150015: READ <= 8'Hd2;
		32'H00150016: READ <= 8'Hc8;
		32'H00150017: READ <= 8'Had;
		32'H00150018: READ <= 8'Haa;
		32'H00150019: READ <= 8'H8f;
		32'H0015001a: READ <= 8'H7a;
		32'H0015001b: READ <= 8'H71;
		32'H0015001c: READ <= 8'H56;
		32'H0015001d: READ <= 8'H7a;
		32'H0015001e: READ <= 8'H75;
		32'H0015001f: READ <= 8'H71;
		32'H00150020: READ <= 8'H65;
		32'H00150021: READ <= 8'H70;
		32'H00150022: READ <= 8'H7d;
		32'H00150023: READ <= 8'H7c;
		32'H00150024: READ <= 8'H42;
		32'H00150025: READ <= 8'He;
		32'H00150026: READ <= 8'H2b;
		32'H00150027: READ <= 8'H2b;
		32'H00150028: READ <= 8'H22;
		32'H00150029: READ <= 8'H29;
		32'H0015002a: READ <= 8'H23;
		32'H0015002b: READ <= 8'H21;
		32'H0015002c: READ <= 8'H23;
		32'H0015002d: READ <= 8'H29;
		32'H0015002e: READ <= 8'H2e;
		32'H0015002f: READ <= 8'H18;
		32'H00150030: READ <= 8'H20;
		32'H00150031: READ <= 8'H38;
		32'H00150032: READ <= 8'H43;
		32'H00150033: READ <= 8'H69;
		32'H00150034: READ <= 8'H77;
		32'H00150035: READ <= 8'H6f;
		32'H00150036: READ <= 8'H5a;
		32'H00150037: READ <= 8'H30;
		32'H00150038: READ <= 8'H3d;
		32'H00150039: READ <= 8'H56;
		32'H0015003a: READ <= 8'H6a;
		32'H0015003b: READ <= 8'H73;
		32'H0015003c: READ <= 8'H72;
		32'H0015003d: READ <= 8'H59;
		32'H0015003e: READ <= 8'H2d;
		32'H0015003f: READ <= 8'H21;
		32'H00150040: READ <= 8'H26;
		32'H00150041: READ <= 8'H33;
		32'H00150042: READ <= 8'H36;
		32'H00150043: READ <= 8'H2a;
		32'H00150044: READ <= 8'H18;
		32'H00150045: READ <= 8'H26;
		32'H00150046: READ <= 8'H3e;
		32'H00150047: READ <= 8'H54;
		32'H00150048: READ <= 8'H79;
		32'H00150049: READ <= 8'H7b;
		32'H0015004a: READ <= 8'H75;
		32'H0015004b: READ <= 8'H7f;
		32'H0015004c: READ <= 8'H8c;
		32'H0015004d: READ <= 8'H8b;
		32'H0015004e: READ <= 8'H88;
		32'H0015004f: READ <= 8'H89;
		32'H00150050: READ <= 8'H8a;
		32'H00150051: READ <= 8'H8b;
		32'H00150052: READ <= 8'H8c;
		32'H00150053: READ <= 8'H8c;
		32'H00150054: READ <= 8'H8c;
		32'H00150055: READ <= 8'H8c;
		32'H00150056: READ <= 8'H8d;
		32'H00150057: READ <= 8'H8c;
		32'H00150058: READ <= 8'H8e;
		32'H00150059: READ <= 8'H8f;
		32'H0015005a: READ <= 8'H8e;
		32'H0015005b: READ <= 8'H90;
		32'H0015005c: READ <= 8'H90;
		32'H0015005d: READ <= 8'H90;
		32'H0015005e: READ <= 8'H90;
		32'H0015005f: READ <= 8'H91;
		32'H00150060: READ <= 8'H90;
		32'H00150061: READ <= 8'H91;
		32'H00150062: READ <= 8'H90;
		32'H00150063: READ <= 8'H8f;
		
		32'H00160000: READ <= 8'H8e;
		32'H00160001: READ <= 8'H90;
		32'H00160002: READ <= 8'H91;
		32'H00160003: READ <= 8'H92;
		32'H00160004: READ <= 8'H95;
		32'H00160005: READ <= 8'H97;
		32'H00160006: READ <= 8'H9b;
		32'H00160007: READ <= 8'Ha0;
		32'H00160008: READ <= 8'Ha3;
		32'H00160009: READ <= 8'Ha8;
		32'H0016000a: READ <= 8'Hac;
		32'H0016000b: READ <= 8'Hae;
		32'H0016000c: READ <= 8'Hb1;
		32'H0016000d: READ <= 8'Hb4;
		32'H0016000e: READ <= 8'Hb8;
		32'H0016000f: READ <= 8'Hbb;
		32'H00160010: READ <= 8'Hbd;
		32'H00160011: READ <= 8'Hbf;
		32'H00160012: READ <= 8'Hc1;
		32'H00160013: READ <= 8'Hc6;
		32'H00160014: READ <= 8'Hcd;
		32'H00160015: READ <= 8'Hcc;
		32'H00160016: READ <= 8'Hb1;
		32'H00160017: READ <= 8'Ha3;
		32'H00160018: READ <= 8'H9f;
		32'H00160019: READ <= 8'H8d;
		32'H0016001a: READ <= 8'H6d;
		32'H0016001b: READ <= 8'H5e;
		32'H0016001c: READ <= 8'H42;
		32'H0016001d: READ <= 8'H68;
		32'H0016001e: READ <= 8'H79;
		32'H0016001f: READ <= 8'H7b;
		32'H00160020: READ <= 8'H5a;
		32'H00160021: READ <= 8'H3c;
		32'H00160022: READ <= 8'H3e;
		32'H00160023: READ <= 8'H35;
		32'H00160024: READ <= 8'H29;
		32'H00160025: READ <= 8'H23;
		32'H00160026: READ <= 8'H1e;
		32'H00160027: READ <= 8'H1b;
		32'H00160028: READ <= 8'H13;
		32'H00160029: READ <= 8'H1d;
		32'H0016002a: READ <= 8'H29;
		32'H0016002b: READ <= 8'H20;
		32'H0016002c: READ <= 8'H3c;
		32'H0016002d: READ <= 8'H40;
		32'H0016002e: READ <= 8'H3f;
		32'H0016002f: READ <= 8'H37;
		32'H00160030: READ <= 8'H5a;
		32'H00160031: READ <= 8'H72;
		32'H00160032: READ <= 8'H72;
		32'H00160033: READ <= 8'H6f;
		32'H00160034: READ <= 8'H7a;
		32'H00160035: READ <= 8'H70;
		32'H00160036: READ <= 8'H63;
		32'H00160037: READ <= 8'H14;
		32'H00160038: READ <= 8'H14;
		32'H00160039: READ <= 8'H20;
		32'H0016003a: READ <= 8'H34;
		32'H0016003b: READ <= 8'H51;
		32'H0016003c: READ <= 8'H62;
		32'H0016003d: READ <= 8'H73;
		32'H0016003e: READ <= 8'H46;
		32'H0016003f: READ <= 8'H38;
		32'H00160040: READ <= 8'H6d;
		32'H00160041: READ <= 8'H3a;
		32'H00160042: READ <= 8'H3c;
		32'H00160043: READ <= 8'H3b;
		32'H00160044: READ <= 8'H2d;
		32'H00160045: READ <= 8'H1f;
		32'H00160046: READ <= 8'H1f;
		32'H00160047: READ <= 8'H37;
		32'H00160048: READ <= 8'H53;
		32'H00160049: READ <= 8'H74;
		32'H0016004a: READ <= 8'H82;
		32'H0016004b: READ <= 8'H77;
		32'H0016004c: READ <= 8'H78;
		32'H0016004d: READ <= 8'H83;
		32'H0016004e: READ <= 8'H8a;
		32'H0016004f: READ <= 8'H88;
		32'H00160050: READ <= 8'H89;
		32'H00160051: READ <= 8'H89;
		32'H00160052: READ <= 8'H8a;
		32'H00160053: READ <= 8'H8a;
		32'H00160054: READ <= 8'H8a;
		32'H00160055: READ <= 8'H8b;
		32'H00160056: READ <= 8'H8c;
		32'H00160057: READ <= 8'H8b;
		32'H00160058: READ <= 8'H8c;
		32'H00160059: READ <= 8'H8d;
		32'H0016005a: READ <= 8'H8e;
		32'H0016005b: READ <= 8'H8e;
		32'H0016005c: READ <= 8'H8f;
		32'H0016005d: READ <= 8'H8e;
		32'H0016005e: READ <= 8'H8f;
		32'H0016005f: READ <= 8'H8f;
		32'H00160060: READ <= 8'H8f;
		32'H00160061: READ <= 8'H8f;
		32'H00160062: READ <= 8'H8e;
		32'H00160063: READ <= 8'H8e;
		
		32'H00170000: READ <= 8'H8e;
		32'H00170001: READ <= 8'H8e;
		32'H00170002: READ <= 8'H8e;
		32'H00170003: READ <= 8'H8f;
		32'H00170004: READ <= 8'H91;
		32'H00170005: READ <= 8'H94;
		32'H00170006: READ <= 8'H98;
		32'H00170007: READ <= 8'H9d;
		32'H00170008: READ <= 8'Ha1;
		32'H00170009: READ <= 8'Ha5;
		32'H0017000a: READ <= 8'Ha9;
		32'H0017000b: READ <= 8'Hac;
		32'H0017000c: READ <= 8'Hae;
		32'H0017000d: READ <= 8'Hb2;
		32'H0017000e: READ <= 8'Hb6;
		32'H0017000f: READ <= 8'Hb9;
		32'H00170010: READ <= 8'Hba;
		32'H00170011: READ <= 8'Hbc;
		32'H00170012: READ <= 8'Hbf;
		32'H00170013: READ <= 8'Hc3;
		32'H00170014: READ <= 8'Hcb;
		32'H00170015: READ <= 8'Hc7;
		32'H00170016: READ <= 8'Haa;
		32'H00170017: READ <= 8'H99;
		32'H00170018: READ <= 8'H9a;
		32'H00170019: READ <= 8'H99;
		32'H0017001a: READ <= 8'H8d;
		32'H0017001b: READ <= 8'H73;
		32'H0017001c: READ <= 8'H53;
		32'H0017001d: READ <= 8'H3f;
		32'H0017001e: READ <= 8'H5e;
		32'H0017001f: READ <= 8'H74;
		32'H00170020: READ <= 8'H55;
		32'H00170021: READ <= 8'H14;
		32'H00170022: READ <= 8'He;
		32'H00170023: READ <= 8'H12;
		32'H00170024: READ <= 8'H14;
		32'H00170025: READ <= 8'H3c;
		32'H00170026: READ <= 8'H5b;
		32'H00170027: READ <= 8'H50;
		32'H00170028: READ <= 8'H45;
		32'H00170029: READ <= 8'H34;
		32'H0017002a: READ <= 8'H1e;
		32'H0017002b: READ <= 8'H3;
		32'H0017002c: READ <= 8'H47;
		32'H0017002d: READ <= 8'H44;
		32'H0017002e: READ <= 8'H32;
		32'H0017002f: READ <= 8'H4c;
		32'H00170030: READ <= 8'H69;
		32'H00170031: READ <= 8'H6a;
		32'H00170032: READ <= 8'H7a;
		32'H00170033: READ <= 8'H78;
		32'H00170034: READ <= 8'H6b;
		32'H00170035: READ <= 8'H72;
		32'H00170036: READ <= 8'H30;
		32'H00170037: READ <= 8'H10;
		32'H00170038: READ <= 8'H10;
		32'H00170039: READ <= 8'H6;
		32'H0017003a: READ <= 8'H2;
		32'H0017003b: READ <= 8'Hd;
		32'H0017003c: READ <= 8'H16;
		32'H0017003d: READ <= 8'H41;
		32'H0017003e: READ <= 8'H50;
		32'H0017003f: READ <= 8'H44;
		32'H00170040: READ <= 8'H82;
		32'H00170041: READ <= 8'H52;
		32'H00170042: READ <= 8'H66;
		32'H00170043: READ <= 8'H65;
		32'H00170044: READ <= 8'H68;
		32'H00170045: READ <= 8'H4d;
		32'H00170046: READ <= 8'H38;
		32'H00170047: READ <= 8'H17;
		32'H00170048: READ <= 8'H21;
		32'H00170049: READ <= 8'H3f;
		32'H0017004a: READ <= 8'H6e;
		32'H0017004b: READ <= 8'H86;
		32'H0017004c: READ <= 8'H7a;
		32'H0017004d: READ <= 8'H74;
		32'H0017004e: READ <= 8'H7e;
		32'H0017004f: READ <= 8'H8a;
		32'H00170050: READ <= 8'H87;
		32'H00170051: READ <= 8'H89;
		32'H00170052: READ <= 8'H89;
		32'H00170053: READ <= 8'H89;
		32'H00170054: READ <= 8'H8a;
		32'H00170055: READ <= 8'H8a;
		32'H00170056: READ <= 8'H8a;
		32'H00170057: READ <= 8'H8a;
		32'H00170058: READ <= 8'H8a;
		32'H00170059: READ <= 8'H8c;
		32'H0017005a: READ <= 8'H8c;
		32'H0017005b: READ <= 8'H8c;
		32'H0017005c: READ <= 8'H8d;
		32'H0017005d: READ <= 8'H8d;
		32'H0017005e: READ <= 8'H8e;
		32'H0017005f: READ <= 8'H8e;
		32'H00170060: READ <= 8'H8d;
		32'H00170061: READ <= 8'H8d;
		32'H00170062: READ <= 8'H8d;
		32'H00170063: READ <= 8'H8c;
		
		32'H00180000: READ <= 8'H8b;
		32'H00180001: READ <= 8'H8b;
		32'H00180002: READ <= 8'H8b;
		32'H00180003: READ <= 8'H8c;
		32'H00180004: READ <= 8'H8e;
		32'H00180005: READ <= 8'H92;
		32'H00180006: READ <= 8'H95;
		32'H00180007: READ <= 8'H9a;
		32'H00180008: READ <= 8'H9f;
		32'H00180009: READ <= 8'Ha2;
		32'H0018000a: READ <= 8'Ha6;
		32'H0018000b: READ <= 8'Ha9;
		32'H0018000c: READ <= 8'Had;
		32'H0018000d: READ <= 8'Hb0;
		32'H0018000e: READ <= 8'Hb3;
		32'H0018000f: READ <= 8'Hb7;
		32'H00180010: READ <= 8'Hb8;
		32'H00180011: READ <= 8'Hba;
		32'H00180012: READ <= 8'Hbc;
		32'H00180013: READ <= 8'Hc2;
		32'H00180014: READ <= 8'Hc5;
		32'H00180015: READ <= 8'Hb3;
		32'H00180016: READ <= 8'H9e;
		32'H00180017: READ <= 8'H98;
		32'H00180018: READ <= 8'H8e;
		32'H00180019: READ <= 8'H8d;
		32'H0018001a: READ <= 8'H93;
		32'H0018001b: READ <= 8'H92;
		32'H0018001c: READ <= 8'H85;
		32'H0018001d: READ <= 8'H52;
		32'H0018001e: READ <= 8'H40;
		32'H0018001f: READ <= 8'H5f;
		32'H00180020: READ <= 8'H54;
		32'H00180021: READ <= 8'H5a;
		32'H00180022: READ <= 8'H71;
		32'H00180023: READ <= 8'H3e;
		32'H00180024: READ <= 8'Ha;
		32'H00180025: READ <= 8'H24;
		32'H00180026: READ <= 8'H5f;
		32'H00180027: READ <= 8'H62;
		32'H00180028: READ <= 8'H59;
		32'H00180029: READ <= 8'H80;
		32'H0018002a: READ <= 8'H5e;
		32'H0018002b: READ <= 8'H54;
		32'H0018002c: READ <= 8'H61;
		32'H0018002d: READ <= 8'H62;
		32'H0018002e: READ <= 8'H5d;
		32'H0018002f: READ <= 8'H4a;
		32'H00180030: READ <= 8'H50;
		32'H00180031: READ <= 8'H76;
		32'H00180032: READ <= 8'H73;
		32'H00180033: READ <= 8'H72;
		32'H00180034: READ <= 8'H6c;
		32'H00180035: READ <= 8'H60;
		32'H00180036: READ <= 8'H3b;
		32'H00180037: READ <= 8'H14;
		32'H00180038: READ <= 8'H6;
		32'H00180039: READ <= 8'H15;
		32'H0018003a: READ <= 8'H2b;
		32'H0018003b: READ <= 8'H14;
		32'H0018003c: READ <= 8'H4;
		32'H0018003d: READ <= 8'H2c;
		32'H0018003e: READ <= 8'H65;
		32'H0018003f: READ <= 8'H82;
		32'H00180040: READ <= 8'H75;
		32'H00180041: READ <= 8'H83;
		32'H00180042: READ <= 8'Hb0;
		32'H00180043: READ <= 8'Ha1;
		32'H00180044: READ <= 8'Hac;
		32'H00180045: READ <= 8'H9c;
		32'H00180046: READ <= 8'H5f;
		32'H00180047: READ <= 8'H4d;
		32'H00180048: READ <= 8'H25;
		32'H00180049: READ <= 8'H2a;
		32'H0018004a: READ <= 8'H36;
		32'H0018004b: READ <= 8'H56;
		32'H0018004c: READ <= 8'H72;
		32'H0018004d: READ <= 8'H84;
		32'H0018004e: READ <= 8'H78;
		32'H0018004f: READ <= 8'H78;
		32'H00180050: READ <= 8'H89;
		32'H00180051: READ <= 8'H87;
		32'H00180052: READ <= 8'H88;
		32'H00180053: READ <= 8'H88;
		32'H00180054: READ <= 8'H89;
		32'H00180055: READ <= 8'H8a;
		32'H00180056: READ <= 8'H8a;
		32'H00180057: READ <= 8'H8a;
		32'H00180058: READ <= 8'H8a;
		32'H00180059: READ <= 8'H8b;
		32'H0018005a: READ <= 8'H8b;
		32'H0018005b: READ <= 8'H8b;
		32'H0018005c: READ <= 8'H8c;
		32'H0018005d: READ <= 8'H8c;
		32'H0018005e: READ <= 8'H8c;
		32'H0018005f: READ <= 8'H8c;
		32'H00180060: READ <= 8'H8b;
		32'H00180061: READ <= 8'H8c;
		32'H00180062: READ <= 8'H8b;
		32'H00180063: READ <= 8'H8b;
		
		32'H00190000: READ <= 8'H89;
		32'H00190001: READ <= 8'H89;
		32'H00190002: READ <= 8'H8a;
		32'H00190003: READ <= 8'H8a;
		32'H00190004: READ <= 8'H8c;
		32'H00190005: READ <= 8'H8f;
		32'H00190006: READ <= 8'H93;
		32'H00190007: READ <= 8'H98;
		32'H00190008: READ <= 8'H9d;
		32'H00190009: READ <= 8'H9f;
		32'H0019000a: READ <= 8'Ha3;
		32'H0019000b: READ <= 8'Ha6;
		32'H0019000c: READ <= 8'Haa;
		32'H0019000d: READ <= 8'Had;
		32'H0019000e: READ <= 8'Hb1;
		32'H0019000f: READ <= 8'Hb3;
		32'H00190010: READ <= 8'Hb6;
		32'H00190011: READ <= 8'Hb8;
		32'H00190012: READ <= 8'Hb9;
		32'H00190013: READ <= 8'Hc1;
		32'H00190014: READ <= 8'Hc9;
		32'H00190015: READ <= 8'Ha7;
		32'H00190016: READ <= 8'H88;
		32'H00190017: READ <= 8'H88;
		32'H00190018: READ <= 8'H8d;
		32'H00190019: READ <= 8'H88;
		32'H0019001a: READ <= 8'H8b;
		32'H0019001b: READ <= 8'H90;
		32'H0019001c: READ <= 8'H96;
		32'H0019001d: READ <= 8'H94;
		32'H0019001e: READ <= 8'H8e;
		32'H0019001f: READ <= 8'H94;
		32'H00190020: READ <= 8'H8c;
		32'H00190021: READ <= 8'H97;
		32'H00190022: READ <= 8'H97;
		32'H00190023: READ <= 8'H81;
		32'H00190024: READ <= 8'H58;
		32'H00190025: READ <= 8'H20;
		32'H00190026: READ <= 8'H42;
		32'H00190027: READ <= 8'H5d;
		32'H00190028: READ <= 8'H79;
		32'H00190029: READ <= 8'H7d;
		32'H0019002a: READ <= 8'H8c;
		32'H0019002b: READ <= 8'H87;
		32'H0019002c: READ <= 8'H70;
		32'H0019002d: READ <= 8'H75;
		32'H0019002e: READ <= 8'H5b;
		32'H0019002f: READ <= 8'H5c;
		32'H00190030: READ <= 8'H5a;
		32'H00190031: READ <= 8'H41;
		32'H00190032: READ <= 8'H78;
		32'H00190033: READ <= 8'H75;
		32'H00190034: READ <= 8'H4d;
		32'H00190035: READ <= 8'H29;
		32'H00190036: READ <= 8'H48;
		32'H00190037: READ <= 8'Hc;
		32'H00190038: READ <= 8'H9;
		32'H00190039: READ <= 8'H26;
		32'H0019003a: READ <= 8'H4a;
		32'H0019003b: READ <= 8'H6f;
		32'H0019003c: READ <= 8'H6;
		32'H0019003d: READ <= 8'Ha;
		32'H0019003e: READ <= 8'H5b;
		32'H0019003f: READ <= 8'Ha3;
		32'H00190040: READ <= 8'H9c;
		32'H00190041: READ <= 8'Haa;
		32'H00190042: READ <= 8'Hb7;
		32'H00190043: READ <= 8'Hc1;
		32'H00190044: READ <= 8'Hc0;
		32'H00190045: READ <= 8'Hbf;
		32'H00190046: READ <= 8'Ha3;
		32'H00190047: READ <= 8'H6f;
		32'H00190048: READ <= 8'H73;
		32'H00190049: READ <= 8'H36;
		32'H0019004a: READ <= 8'H30;
		32'H0019004b: READ <= 8'H51;
		32'H0019004c: READ <= 8'H3a;
		32'H0019004d: READ <= 8'H41;
		32'H0019004e: READ <= 8'H74;
		32'H0019004f: READ <= 8'H8d;
		32'H00190050: READ <= 8'H7b;
		32'H00190051: READ <= 8'H88;
		32'H00190052: READ <= 8'H88;
		32'H00190053: READ <= 8'H88;
		32'H00190054: READ <= 8'H88;
		32'H00190055: READ <= 8'H88;
		32'H00190056: READ <= 8'H89;
		32'H00190057: READ <= 8'H89;
		32'H00190058: READ <= 8'H89;
		32'H00190059: READ <= 8'H89;
		32'H0019005a: READ <= 8'H89;
		32'H0019005b: READ <= 8'H8a;
		32'H0019005c: READ <= 8'H8a;
		32'H0019005d: READ <= 8'H8a;
		32'H0019005e: READ <= 8'H8a;
		32'H0019005f: READ <= 8'H8a;
		32'H00190060: READ <= 8'H8b;
		32'H00190061: READ <= 8'H8b;
		32'H00190062: READ <= 8'H8a;
		32'H00190063: READ <= 8'H8a;
		
		32'H001a0000: READ <= 8'H87;
		32'H001a0001: READ <= 8'H87;
		32'H001a0002: READ <= 8'H89;
		32'H001a0003: READ <= 8'H89;
		32'H001a0004: READ <= 8'H8a;
		32'H001a0005: READ <= 8'H8c;
		32'H001a0006: READ <= 8'H91;
		32'H001a0007: READ <= 8'H95;
		32'H001a0008: READ <= 8'H99;
		32'H001a0009: READ <= 8'H9d;
		32'H001a000a: READ <= 8'H9f;
		32'H001a000b: READ <= 8'Ha3;
		32'H001a000c: READ <= 8'Ha7;
		32'H001a000d: READ <= 8'Hab;
		32'H001a000e: READ <= 8'Haf;
		32'H001a000f: READ <= 8'Hb2;
		32'H001a0010: READ <= 8'Hb4;
		32'H001a0011: READ <= 8'Hb5;
		32'H001a0012: READ <= 8'Hb7;
		32'H001a0013: READ <= 8'Hc1;
		32'H001a0014: READ <= 8'Hc3;
		32'H001a0015: READ <= 8'H99;
		32'H001a0016: READ <= 8'H80;
		32'H001a0017: READ <= 8'H85;
		32'H001a0018: READ <= 8'H7f;
		32'H001a0019: READ <= 8'H85;
		32'H001a001a: READ <= 8'H86;
		32'H001a001b: READ <= 8'H86;
		32'H001a001c: READ <= 8'H8e;
		32'H001a001d: READ <= 8'H8f;
		32'H001a001e: READ <= 8'H90;
		32'H001a001f: READ <= 8'H8a;
		32'H001a0020: READ <= 8'H95;
		32'H001a0021: READ <= 8'H98;
		32'H001a0022: READ <= 8'H88;
		32'H001a0023: READ <= 8'H73;
		32'H001a0024: READ <= 8'H79;
		32'H001a0025: READ <= 8'H4d;
		32'H001a0026: READ <= 8'H5a;
		32'H001a0027: READ <= 8'H6b;
		32'H001a0028: READ <= 8'H81;
		32'H001a0029: READ <= 8'H7c;
		32'H001a002a: READ <= 8'H71;
		32'H001a002b: READ <= 8'H6f;
		32'H001a002c: READ <= 8'H6d;
		32'H001a002d: READ <= 8'H7d;
		32'H001a002e: READ <= 8'H79;
		32'H001a002f: READ <= 8'H66;
		32'H001a0030: READ <= 8'H55;
		32'H001a0031: READ <= 8'H3c;
		32'H001a0032: READ <= 8'H4e;
		32'H001a0033: READ <= 8'H47;
		32'H001a0034: READ <= 8'H10;
		32'H001a0035: READ <= 8'H32;
		32'H001a0036: READ <= 8'H43;
		32'H001a0037: READ <= 8'Hd;
		32'H001a0038: READ <= 8'H8;
		32'H001a0039: READ <= 8'H34;
		32'H001a003a: READ <= 8'H46;
		32'H001a003b: READ <= 8'H8f;
		32'H001a003c: READ <= 8'H35;
		32'H001a003d: READ <= 8'H0;
		32'H001a003e: READ <= 8'H49;
		32'H001a003f: READ <= 8'Hab;
		32'H001a0040: READ <= 8'Hb8;
		32'H001a0041: READ <= 8'Hbb;
		32'H001a0042: READ <= 8'Hba;
		32'H001a0043: READ <= 8'Hc1;
		32'H001a0044: READ <= 8'Hb7;
		32'H001a0045: READ <= 8'Hbd;
		32'H001a0046: READ <= 8'Hc5;
		32'H001a0047: READ <= 8'H93;
		32'H001a0048: READ <= 8'H87;
		32'H001a0049: READ <= 8'H80;
		32'H001a004a: READ <= 8'H6c;
		32'H001a004b: READ <= 8'H49;
		32'H001a004c: READ <= 8'H43;
		32'H001a004d: READ <= 8'H2b;
		32'H001a004e: READ <= 8'H28;
		32'H001a004f: READ <= 8'H4b;
		32'H001a0050: READ <= 8'H80;
		32'H001a0051: READ <= 8'H92;
		32'H001a0052: READ <= 8'H89;
		32'H001a0053: READ <= 8'H87;
		32'H001a0054: READ <= 8'H87;
		32'H001a0055: READ <= 8'H88;
		32'H001a0056: READ <= 8'H88;
		32'H001a0057: READ <= 8'H88;
		32'H001a0058: READ <= 8'H88;
		32'H001a0059: READ <= 8'H88;
		32'H001a005a: READ <= 8'H88;
		32'H001a005b: READ <= 8'H88;
		32'H001a005c: READ <= 8'H89;
		32'H001a005d: READ <= 8'H88;
		32'H001a005e: READ <= 8'H89;
		32'H001a005f: READ <= 8'H88;
		32'H001a0060: READ <= 8'H89;
		32'H001a0061: READ <= 8'H8a;
		32'H001a0062: READ <= 8'H8a;
		32'H001a0063: READ <= 8'H89;
		
		32'H001b0000: READ <= 8'H85;
		32'H001b0001: READ <= 8'H86;
		32'H001b0002: READ <= 8'H87;
		32'H001b0003: READ <= 8'H88;
		32'H001b0004: READ <= 8'H88;
		32'H001b0005: READ <= 8'H8b;
		32'H001b0006: READ <= 8'H8d;
		32'H001b0007: READ <= 8'H91;
		32'H001b0008: READ <= 8'H95;
		32'H001b0009: READ <= 8'H9a;
		32'H001b000a: READ <= 8'H9d;
		32'H001b000b: READ <= 8'Ha0;
		32'H001b000c: READ <= 8'Ha5;
		32'H001b000d: READ <= 8'Ha8;
		32'H001b000e: READ <= 8'Hac;
		32'H001b000f: READ <= 8'Hb0;
		32'H001b0010: READ <= 8'Hb1;
		32'H001b0011: READ <= 8'Hb3;
		32'H001b0012: READ <= 8'Hb6;
		32'H001b0013: READ <= 8'Hc0;
		32'H001b0014: READ <= 8'Hc2;
		32'H001b0015: READ <= 8'H92;
		32'H001b0016: READ <= 8'H89;
		32'H001b0017: READ <= 8'H89;
		32'H001b0018: READ <= 8'H76;
		32'H001b0019: READ <= 8'H7b;
		32'H001b001a: READ <= 8'H78;
		32'H001b001b: READ <= 8'H7b;
		32'H001b001c: READ <= 8'H8d;
		32'H001b001d: READ <= 8'H8a;
		32'H001b001e: READ <= 8'H8d;
		32'H001b001f: READ <= 8'H80;
		32'H001b0020: READ <= 8'H76;
		32'H001b0021: READ <= 8'H7a;
		32'H001b0022: READ <= 8'H80;
		32'H001b0023: READ <= 8'H72;
		32'H001b0024: READ <= 8'H75;
		32'H001b0025: READ <= 8'H34;
		32'H001b0026: READ <= 8'H49;
		32'H001b0027: READ <= 8'H6b;
		32'H001b0028: READ <= 8'H52;
		32'H001b0029: READ <= 8'H55;
		32'H001b002a: READ <= 8'H68;
		32'H001b002b: READ <= 8'H70;
		32'H001b002c: READ <= 8'H6f;
		32'H001b002d: READ <= 8'H61;
		32'H001b002e: READ <= 8'H74;
		32'H001b002f: READ <= 8'H6f;
		32'H001b0030: READ <= 8'H4e;
		32'H001b0031: READ <= 8'H4c;
		32'H001b0032: READ <= 8'H24;
		32'H001b0033: READ <= 8'H7;
		32'H001b0034: READ <= 8'H1a;
		32'H001b0035: READ <= 8'H43;
		32'H001b0036: READ <= 8'H49;
		32'H001b0037: READ <= 8'H9;
		32'H001b0038: READ <= 8'H6;
		32'H001b0039: READ <= 8'H18;
		32'H001b003a: READ <= 8'H62;
		32'H001b003b: READ <= 8'H94;
		32'H001b003c: READ <= 8'Haf;
		32'H001b003d: READ <= 8'H5;
		32'H001b003e: READ <= 8'H31;
		32'H001b003f: READ <= 8'Ha3;
		32'H001b0040: READ <= 8'H9d;
		32'H001b0041: READ <= 8'Hb2;
		32'H001b0042: READ <= 8'Hb6;
		32'H001b0043: READ <= 8'Hba;
		32'H001b0044: READ <= 8'Hbf;
		32'H001b0045: READ <= 8'Hc1;
		32'H001b0046: READ <= 8'Hbf;
		32'H001b0047: READ <= 8'Hb3;
		32'H001b0048: READ <= 8'H84;
		32'H001b0049: READ <= 8'H94;
		32'H001b004a: READ <= 8'H93;
		32'H001b004b: READ <= 8'H8d;
		32'H001b004c: READ <= 8'H74;
		32'H001b004d: READ <= 8'H84;
		32'H001b004e: READ <= 8'H51;
		32'H001b004f: READ <= 8'H38;
		32'H001b0050: READ <= 8'H32;
		32'H001b0051: READ <= 8'H5b;
		32'H001b0052: READ <= 8'H7d;
		32'H001b0053: READ <= 8'H87;
		32'H001b0054: READ <= 8'H86;
		32'H001b0055: READ <= 8'H87;
		32'H001b0056: READ <= 8'H87;
		32'H001b0057: READ <= 8'H87;
		32'H001b0058: READ <= 8'H88;
		32'H001b0059: READ <= 8'H87;
		32'H001b005a: READ <= 8'H87;
		32'H001b005b: READ <= 8'H88;
		32'H001b005c: READ <= 8'H88;
		32'H001b005d: READ <= 8'H87;
		32'H001b005e: READ <= 8'H88;
		32'H001b005f: READ <= 8'H88;
		32'H001b0060: READ <= 8'H88;
		32'H001b0061: READ <= 8'H88;
		32'H001b0062: READ <= 8'H89;
		32'H001b0063: READ <= 8'H89;
		
		32'H001c0000: READ <= 8'H83;
		32'H001c0001: READ <= 8'H84;
		32'H001c0002: READ <= 8'H85;
		32'H001c0003: READ <= 8'H87;
		32'H001c0004: READ <= 8'H87;
		32'H001c0005: READ <= 8'H89;
		32'H001c0006: READ <= 8'H8c;
		32'H001c0007: READ <= 8'H8f;
		32'H001c0008: READ <= 8'H93;
		32'H001c0009: READ <= 8'H97;
		32'H001c000a: READ <= 8'H9b;
		32'H001c000b: READ <= 8'H9e;
		32'H001c000c: READ <= 8'Ha3;
		32'H001c000d: READ <= 8'Ha5;
		32'H001c000e: READ <= 8'Ha9;
		32'H001c000f: READ <= 8'Hac;
		32'H001c0010: READ <= 8'Haf;
		32'H001c0011: READ <= 8'Hb0;
		32'H001c0012: READ <= 8'Hb3;
		32'H001c0013: READ <= 8'Hbe;
		32'H001c0014: READ <= 8'Hc5;
		32'H001c0015: READ <= 8'Ha0;
		32'H001c0016: READ <= 8'H91;
		32'H001c0017: READ <= 8'H78;
		32'H001c0018: READ <= 8'H7e;
		32'H001c0019: READ <= 8'H74;
		32'H001c001a: READ <= 8'H72;
		32'H001c001b: READ <= 8'H82;
		32'H001c001c: READ <= 8'H77;
		32'H001c001d: READ <= 8'H8b;
		32'H001c001e: READ <= 8'H7b;
		32'H001c001f: READ <= 8'H85;
		32'H001c0020: READ <= 8'H76;
		32'H001c0021: READ <= 8'H80;
		32'H001c0022: READ <= 8'H62;
		32'H001c0023: READ <= 8'H56;
		32'H001c0024: READ <= 8'H16;
		32'H001c0025: READ <= 8'H14;
		32'H001c0026: READ <= 8'H45;
		32'H001c0027: READ <= 8'H6b;
		32'H001c0028: READ <= 8'H65;
		32'H001c0029: READ <= 8'H68;
		32'H001c002a: READ <= 8'H65;
		32'H001c002b: READ <= 8'H61;
		32'H001c002c: READ <= 8'H5f;
		32'H001c002d: READ <= 8'H69;
		32'H001c002e: READ <= 8'H72;
		32'H001c002f: READ <= 8'H8a;
		32'H001c0030: READ <= 8'H5d;
		32'H001c0031: READ <= 8'H4e;
		32'H001c0032: READ <= 8'H22;
		32'H001c0033: READ <= 8'H1;
		32'H001c0034: READ <= 8'H22;
		32'H001c0035: READ <= 8'H53;
		32'H001c0036: READ <= 8'H49;
		32'H001c0037: READ <= 8'H9;
		32'H001c0038: READ <= 8'H6;
		32'H001c0039: READ <= 8'H1b;
		32'H001c003a: READ <= 8'H67;
		32'H001c003b: READ <= 8'H85;
		32'H001c003c: READ <= 8'Hb4;
		32'H001c003d: READ <= 8'H45;
		32'H001c003e: READ <= 8'H1b;
		32'H001c003f: READ <= 8'H9f;
		32'H001c0040: READ <= 8'Hb6;
		32'H001c0041: READ <= 8'Ha8;
		32'H001c0042: READ <= 8'Hb1;
		32'H001c0043: READ <= 8'Hb4;
		32'H001c0044: READ <= 8'Hb7;
		32'H001c0045: READ <= 8'Hbf;
		32'H001c0046: READ <= 8'Hc2;
		32'H001c0047: READ <= 8'Hb9;
		32'H001c0048: READ <= 8'H8b;
		32'H001c0049: READ <= 8'H65;
		32'H001c004a: READ <= 8'H8c;
		32'H001c004b: READ <= 8'Ha4;
		32'H001c004c: READ <= 8'Ha0;
		32'H001c004d: READ <= 8'Ha0;
		32'H001c004e: READ <= 8'H9a;
		32'H001c004f: READ <= 8'H54;
		32'H001c0050: READ <= 8'H49;
		32'H001c0051: READ <= 8'H47;
		32'H001c0052: READ <= 8'H40;
		32'H001c0053: READ <= 8'H58;
		32'H001c0054: READ <= 8'H85;
		32'H001c0055: READ <= 8'H87;
		32'H001c0056: READ <= 8'H86;
		32'H001c0057: READ <= 8'H86;
		32'H001c0058: READ <= 8'H86;
		32'H001c0059: READ <= 8'H86;
		32'H001c005a: READ <= 8'H86;
		32'H001c005b: READ <= 8'H87;
		32'H001c005c: READ <= 8'H87;
		32'H001c005d: READ <= 8'H86;
		32'H001c005e: READ <= 8'H88;
		32'H001c005f: READ <= 8'H87;
		32'H001c0060: READ <= 8'H87;
		32'H001c0061: READ <= 8'H88;
		32'H001c0062: READ <= 8'H88;
		32'H001c0063: READ <= 8'H89;
		
		32'H001d0000: READ <= 8'H83;
		32'H001d0001: READ <= 8'H83;
		32'H001d0002: READ <= 8'H84;
		32'H001d0003: READ <= 8'H84;
		32'H001d0004: READ <= 8'H85;
		32'H001d0005: READ <= 8'H87;
		32'H001d0006: READ <= 8'H89;
		32'H001d0007: READ <= 8'H8b;
		32'H001d0008: READ <= 8'H90;
		32'H001d0009: READ <= 8'H93;
		32'H001d000a: READ <= 8'H98;
		32'H001d000b: READ <= 8'H9b;
		32'H001d000c: READ <= 8'Ha0;
		32'H001d000d: READ <= 8'Ha3;
		32'H001d000e: READ <= 8'Ha6;
		32'H001d000f: READ <= 8'Ha8;
		32'H001d0010: READ <= 8'Hac;
		32'H001d0011: READ <= 8'Hae;
		32'H001d0012: READ <= 8'Hb2;
		32'H001d0013: READ <= 8'Hbb;
		32'H001d0014: READ <= 8'Hc1;
		32'H001d0015: READ <= 8'H9e;
		32'H001d0016: READ <= 8'H82;
		32'H001d0017: READ <= 8'H84;
		32'H001d0018: READ <= 8'H79;
		32'H001d0019: READ <= 8'H74;
		32'H001d001a: READ <= 8'H73;
		32'H001d001b: READ <= 8'H7d;
		32'H001d001c: READ <= 8'H7b;
		32'H001d001d: READ <= 8'H8c;
		32'H001d001e: READ <= 8'H84;
		32'H001d001f: READ <= 8'H7d;
		32'H001d0020: READ <= 8'H70;
		32'H001d0021: READ <= 8'H6a;
		32'H001d0022: READ <= 8'H55;
		32'H001d0023: READ <= 8'H13;
		32'H001d0024: READ <= 8'H8;
		32'H001d0025: READ <= 8'H1b;
		32'H001d0026: READ <= 8'H44;
		32'H001d0027: READ <= 8'H5a;
		32'H001d0028: READ <= 8'H4d;
		32'H001d0029: READ <= 8'H51;
		32'H001d002a: READ <= 8'H59;
		32'H001d002b: READ <= 8'H5e;
		32'H001d002c: READ <= 8'H82;
		32'H001d002d: READ <= 8'H69;
		32'H001d002e: READ <= 8'H5c;
		32'H001d002f: READ <= 8'H5f;
		32'H001d0030: READ <= 8'H65;
		32'H001d0031: READ <= 8'H50;
		32'H001d0032: READ <= 8'H2b;
		32'H001d0033: READ <= 8'H15;
		32'H001d0034: READ <= 8'H32;
		32'H001d0035: READ <= 8'H61;
		32'H001d0036: READ <= 8'H43;
		32'H001d0037: READ <= 8'Hc;
		32'H001d0038: READ <= 8'Ha;
		32'H001d0039: READ <= 8'H1b;
		32'H001d003a: READ <= 8'H63;
		32'H001d003b: READ <= 8'H8c;
		32'H001d003c: READ <= 8'Ha0;
		32'H001d003d: READ <= 8'H6e;
		32'H001d003e: READ <= 8'Hb;
		32'H001d003f: READ <= 8'H76;
		32'H001d0040: READ <= 8'Ha4;
		32'H001d0041: READ <= 8'Haa;
		32'H001d0042: READ <= 8'Hac;
		32'H001d0043: READ <= 8'Hac;
		32'H001d0044: READ <= 8'Hb7;
		32'H001d0045: READ <= 8'Hba;
		32'H001d0046: READ <= 8'Hc0;
		32'H001d0047: READ <= 8'Hb9;
		32'H001d0048: READ <= 8'H97;
		32'H001d0049: READ <= 8'H4e;
		32'H001d004a: READ <= 8'H4f;
		32'H001d004b: READ <= 8'Ha4;
		32'H001d004c: READ <= 8'Hb0;
		32'H001d004d: READ <= 8'Ha6;
		32'H001d004e: READ <= 8'Ha9;
		32'H001d004f: READ <= 8'H99;
		32'H001d0050: READ <= 8'H7f;
		32'H001d0051: READ <= 8'H92;
		32'H001d0052: READ <= 8'H64;
		32'H001d0053: READ <= 8'H4c;
		32'H001d0054: READ <= 8'H5a;
		32'H001d0055: READ <= 8'H85;
		32'H001d0056: READ <= 8'H87;
		32'H001d0057: READ <= 8'H86;
		32'H001d0058: READ <= 8'H86;
		32'H001d0059: READ <= 8'H86;
		32'H001d005a: READ <= 8'H86;
		32'H001d005b: READ <= 8'H86;
		32'H001d005c: READ <= 8'H86;
		32'H001d005d: READ <= 8'H86;
		32'H001d005e: READ <= 8'H87;
		32'H001d005f: READ <= 8'H87;
		32'H001d0060: READ <= 8'H87;
		32'H001d0061: READ <= 8'H88;
		32'H001d0062: READ <= 8'H88;
		32'H001d0063: READ <= 8'H88;
		
		32'H001e0000: READ <= 8'H82;
		32'H001e0001: READ <= 8'H82;
		32'H001e0002: READ <= 8'H82;
		32'H001e0003: READ <= 8'H83;
		32'H001e0004: READ <= 8'H84;
		32'H001e0005: READ <= 8'H85;
		32'H001e0006: READ <= 8'H87;
		32'H001e0007: READ <= 8'H89;
		32'H001e0008: READ <= 8'H8d;
		32'H001e0009: READ <= 8'H90;
		32'H001e000a: READ <= 8'H95;
		32'H001e000b: READ <= 8'H99;
		32'H001e000c: READ <= 8'H9c;
		32'H001e000d: READ <= 8'H9f;
		32'H001e000e: READ <= 8'Ha2;
		32'H001e000f: READ <= 8'Ha5;
		32'H001e0010: READ <= 8'Ha9;
		32'H001e0011: READ <= 8'Hab;
		32'H001e0012: READ <= 8'Hac;
		32'H001e0013: READ <= 8'Hbb;
		32'H001e0014: READ <= 8'Hc9;
		32'H001e0015: READ <= 8'H99;
		32'H001e0016: READ <= 8'H83;
		32'H001e0017: READ <= 8'H78;
		32'H001e0018: READ <= 8'H71;
		32'H001e0019: READ <= 8'H6b;
		32'H001e001a: READ <= 8'H72;
		32'H001e001b: READ <= 8'H74;
		32'H001e001c: READ <= 8'H74;
		32'H001e001d: READ <= 8'H81;
		32'H001e001e: READ <= 8'H7d;
		32'H001e001f: READ <= 8'H75;
		32'H001e0020: READ <= 8'H6f;
		32'H001e0021: READ <= 8'H63;
		32'H001e0022: READ <= 8'H3b;
		32'H001e0023: READ <= 8'H20;
		32'H001e0024: READ <= 8'H13;
		32'H001e0025: READ <= 8'H6;
		32'H001e0026: READ <= 8'H3c;
		32'H001e0027: READ <= 8'H4f;
		32'H001e0028: READ <= 8'H51;
		32'H001e0029: READ <= 8'H4c;
		32'H001e002a: READ <= 8'H6c;
		32'H001e002b: READ <= 8'H6d;
		32'H001e002c: READ <= 8'H72;
		32'H001e002d: READ <= 8'H7d;
		32'H001e002e: READ <= 8'H6e;
		32'H001e002f: READ <= 8'H7c;
		32'H001e0030: READ <= 8'H4a;
		32'H001e0031: READ <= 8'H41;
		32'H001e0032: READ <= 8'H19;
		32'H001e0033: READ <= 8'H2b;
		32'H001e0034: READ <= 8'H31;
		32'H001e0035: READ <= 8'H60;
		32'H001e0036: READ <= 8'H3c;
		32'H001e0037: READ <= 8'H8;
		32'H001e0038: READ <= 8'H6;
		32'H001e0039: READ <= 8'H1a;
		32'H001e003a: READ <= 8'H63;
		32'H001e003b: READ <= 8'H82;
		32'H001e003c: READ <= 8'H8d;
		32'H001e003d: READ <= 8'H7a;
		32'H001e003e: READ <= 8'H0;
		32'H001e003f: READ <= 8'H63;
		32'H001e0040: READ <= 8'Ha1;
		32'H001e0041: READ <= 8'H9d;
		32'H001e0042: READ <= 8'H9b;
		32'H001e0043: READ <= 8'Ha5;
		32'H001e0044: READ <= 8'Haa;
		32'H001e0045: READ <= 8'Had;
		32'H001e0046: READ <= 8'Hb7;
		32'H001e0047: READ <= 8'Hb5;
		32'H001e0048: READ <= 8'H98;
		32'H001e0049: READ <= 8'H4f;
		32'H001e004a: READ <= 8'H39;
		32'H001e004b: READ <= 8'H69;
		32'H001e004c: READ <= 8'Ha8;
		32'H001e004d: READ <= 8'Hb4;
		32'H001e004e: READ <= 8'Had;
		32'H001e004f: READ <= 8'Ha0;
		32'H001e0050: READ <= 8'H97;
		32'H001e0051: READ <= 8'H95;
		32'H001e0052: READ <= 8'H92;
		32'H001e0053: READ <= 8'H6f;
		32'H001e0054: READ <= 8'H5a;
		32'H001e0055: READ <= 8'H67;
		32'H001e0056: READ <= 8'H89;
		32'H001e0057: READ <= 8'H85;
		32'H001e0058: READ <= 8'H85;
		32'H001e0059: READ <= 8'H85;
		32'H001e005a: READ <= 8'H84;
		32'H001e005b: READ <= 8'H85;
		32'H001e005c: READ <= 8'H85;
		32'H001e005d: READ <= 8'H86;
		32'H001e005e: READ <= 8'H86;
		32'H001e005f: READ <= 8'H87;
		32'H001e0060: READ <= 8'H87;
		32'H001e0061: READ <= 8'H87;
		32'H001e0062: READ <= 8'H88;
		32'H001e0063: READ <= 8'H88;
		
		32'H001f0000: READ <= 8'H81;
		32'H001f0001: READ <= 8'H81;
		32'H001f0002: READ <= 8'H81;
		32'H001f0003: READ <= 8'H81;
		32'H001f0004: READ <= 8'H82;
		32'H001f0005: READ <= 8'H83;
		32'H001f0006: READ <= 8'H84;
		32'H001f0007: READ <= 8'H86;
		32'H001f0008: READ <= 8'H8a;
		32'H001f0009: READ <= 8'H8e;
		32'H001f000a: READ <= 8'H91;
		32'H001f000b: READ <= 8'H95;
		32'H001f000c: READ <= 8'H99;
		32'H001f000d: READ <= 8'H9c;
		32'H001f000e: READ <= 8'H9f;
		32'H001f000f: READ <= 8'Ha1;
		32'H001f0010: READ <= 8'Ha5;
		32'H001f0011: READ <= 8'Ha8;
		32'H001f0012: READ <= 8'Haa;
		32'H001f0013: READ <= 8'Hb1;
		32'H001f0014: READ <= 8'Hc5;
		32'H001f0015: READ <= 8'Ha0;
		32'H001f0016: READ <= 8'H80;
		32'H001f0017: READ <= 8'H71;
		32'H001f0018: READ <= 8'H6a;
		32'H001f0019: READ <= 8'H77;
		32'H001f001a: READ <= 8'H77;
		32'H001f001b: READ <= 8'H77;
		32'H001f001c: READ <= 8'H6d;
		32'H001f001d: READ <= 8'H6f;
		32'H001f001e: READ <= 8'H76;
		32'H001f001f: READ <= 8'H74;
		32'H001f0020: READ <= 8'H59;
		32'H001f0021: READ <= 8'H51;
		32'H001f0022: READ <= 8'H35;
		32'H001f0023: READ <= 8'H33;
		32'H001f0024: READ <= 8'H9;
		32'H001f0025: READ <= 8'H1;
		32'H001f0026: READ <= 8'H9;
		32'H001f0027: READ <= 8'H4b;
		32'H001f0028: READ <= 8'H45;
		32'H001f0029: READ <= 8'H56;
		32'H001f002a: READ <= 8'H50;
		32'H001f002b: READ <= 8'H60;
		32'H001f002c: READ <= 8'H67;
		32'H001f002d: READ <= 8'H58;
		32'H001f002e: READ <= 8'H64;
		32'H001f002f: READ <= 8'H5a;
		32'H001f0030: READ <= 8'H63;
		32'H001f0031: READ <= 8'H51;
		32'H001f0032: READ <= 8'H1b;
		32'H001f0033: READ <= 8'H36;
		32'H001f0034: READ <= 8'H34;
		32'H001f0035: READ <= 8'H66;
		32'H001f0036: READ <= 8'H2e;
		32'H001f0037: READ <= 8'H5;
		32'H001f0038: READ <= 8'H6;
		32'H001f0039: READ <= 8'H21;
		32'H001f003a: READ <= 8'H6c;
		32'H001f003b: READ <= 8'H82;
		32'H001f003c: READ <= 8'H90;
		32'H001f003d: READ <= 8'H7e;
		32'H001f003e: READ <= 8'H1;
		32'H001f003f: READ <= 8'H28;
		32'H001f0040: READ <= 8'H9a;
		32'H001f0041: READ <= 8'Ha7;
		32'H001f0042: READ <= 8'H9f;
		32'H001f0043: READ <= 8'H9d;
		32'H001f0044: READ <= 8'Hab;
		32'H001f0045: READ <= 8'Ha7;
		32'H001f0046: READ <= 8'Haa;
		32'H001f0047: READ <= 8'Ha8;
		32'H001f0048: READ <= 8'H8f;
		32'H001f0049: READ <= 8'H54;
		32'H001f004a: READ <= 8'H5e;
		32'H001f004b: READ <= 8'H4d;
		32'H001f004c: READ <= 8'H6b;
		32'H001f004d: READ <= 8'Ha0;
		32'H001f004e: READ <= 8'Ha6;
		32'H001f004f: READ <= 8'Ha7;
		32'H001f0050: READ <= 8'H8f;
		32'H001f0051: READ <= 8'Ha3;
		32'H001f0052: READ <= 8'Ha4;
		32'H001f0053: READ <= 8'H91;
		32'H001f0054: READ <= 8'H73;
		32'H001f0055: READ <= 8'H63;
		32'H001f0056: READ <= 8'H6f;
		32'H001f0057: READ <= 8'H86;
		32'H001f0058: READ <= 8'H86;
		32'H001f0059: READ <= 8'H84;
		32'H001f005a: READ <= 8'H84;
		32'H001f005b: READ <= 8'H85;
		32'H001f005c: READ <= 8'H85;
		32'H001f005d: READ <= 8'H85;
		32'H001f005e: READ <= 8'H86;
		32'H001f005f: READ <= 8'H86;
		32'H001f0060: READ <= 8'H88;
		32'H001f0061: READ <= 8'H87;
		32'H001f0062: READ <= 8'H88;
		32'H001f0063: READ <= 8'H88;
		
		32'H00200000: READ <= 8'H7f;
		32'H00200001: READ <= 8'H80;
		32'H00200002: READ <= 8'H80;
		32'H00200003: READ <= 8'H80;
		32'H00200004: READ <= 8'H80;
		32'H00200005: READ <= 8'H81;
		32'H00200006: READ <= 8'H82;
		32'H00200007: READ <= 8'H84;
		32'H00200008: READ <= 8'H87;
		32'H00200009: READ <= 8'H89;
		32'H0020000a: READ <= 8'H8d;
		32'H0020000b: READ <= 8'H92;
		32'H0020000c: READ <= 8'H95;
		32'H0020000d: READ <= 8'H98;
		32'H0020000e: READ <= 8'H9c;
		32'H0020000f: READ <= 8'H9e;
		32'H00200010: READ <= 8'Ha2;
		32'H00200011: READ <= 8'Ha4;
		32'H00200012: READ <= 8'Ha6;
		32'H00200013: READ <= 8'Hba;
		32'H00200014: READ <= 8'Hcf;
		32'H00200015: READ <= 8'Ha2;
		32'H00200016: READ <= 8'H7d;
		32'H00200017: READ <= 8'H6b;
		32'H00200018: READ <= 8'H6e;
		32'H00200019: READ <= 8'H6d;
		32'H0020001a: READ <= 8'H74;
		32'H0020001b: READ <= 8'H6b;
		32'H0020001c: READ <= 8'H76;
		32'H0020001d: READ <= 8'H7e;
		32'H0020001e: READ <= 8'H6a;
		32'H0020001f: READ <= 8'H66;
		32'H00200020: READ <= 8'H69;
		32'H00200021: READ <= 8'H54;
		32'H00200022: READ <= 8'H29;
		32'H00200023: READ <= 8'H2d;
		32'H00200024: READ <= 8'H7;
		32'H00200025: READ <= 8'H7;
		32'H00200026: READ <= 8'H2;
		32'H00200027: READ <= 8'H3f;
		32'H00200028: READ <= 8'H3f;
		32'H00200029: READ <= 8'H51;
		32'H0020002a: READ <= 8'H59;
		32'H0020002b: READ <= 8'H4e;
		32'H0020002c: READ <= 8'H6a;
		32'H0020002d: READ <= 8'H67;
		32'H0020002e: READ <= 8'H65;
		32'H0020002f: READ <= 8'H58;
		32'H00200030: READ <= 8'H46;
		32'H00200031: READ <= 8'H55;
		32'H00200032: READ <= 8'H1a;
		32'H00200033: READ <= 8'H40;
		32'H00200034: READ <= 8'H41;
		32'H00200035: READ <= 8'H67;
		32'H00200036: READ <= 8'H1f;
		32'H00200037: READ <= 8'H3;
		32'H00200038: READ <= 8'H5;
		32'H00200039: READ <= 8'H28;
		32'H0020003a: READ <= 8'H74;
		32'H0020003b: READ <= 8'H7a;
		32'H0020003c: READ <= 8'H95;
		32'H0020003d: READ <= 8'H93;
		32'H0020003e: READ <= 8'H2;
		32'H0020003f: READ <= 8'H3;
		32'H00200040: READ <= 8'H76;
		32'H00200041: READ <= 8'H9a;
		32'H00200042: READ <= 8'Ha2;
		32'H00200043: READ <= 8'Ha5;
		32'H00200044: READ <= 8'Ha1;
		32'H00200045: READ <= 8'H9f;
		32'H00200046: READ <= 8'H99;
		32'H00200047: READ <= 8'H9a;
		32'H00200048: READ <= 8'H81;
		32'H00200049: READ <= 8'H71;
		32'H0020004a: READ <= 8'H72;
		32'H0020004b: READ <= 8'H70;
		32'H0020004c: READ <= 8'H48;
		32'H0020004d: READ <= 8'H77;
		32'H0020004e: READ <= 8'H8c;
		32'H0020004f: READ <= 8'Hac;
		32'H00200050: READ <= 8'H9d;
		32'H00200051: READ <= 8'H95;
		32'H00200052: READ <= 8'Ha8;
		32'H00200053: READ <= 8'Hab;
		32'H00200054: READ <= 8'H94;
		32'H00200055: READ <= 8'H73;
		32'H00200056: READ <= 8'H68;
		32'H00200057: READ <= 8'H72;
		32'H00200058: READ <= 8'H80;
		32'H00200059: READ <= 8'H87;
		32'H0020005a: READ <= 8'H84;
		32'H0020005b: READ <= 8'H85;
		32'H0020005c: READ <= 8'H85;
		32'H0020005d: READ <= 8'H86;
		32'H0020005e: READ <= 8'H86;
		32'H0020005f: READ <= 8'H87;
		32'H00200060: READ <= 8'H87;
		32'H00200061: READ <= 8'H88;
		32'H00200062: READ <= 8'H88;
		32'H00200063: READ <= 8'H88;
		
		32'H00210000: READ <= 8'H7e;
		32'H00210001: READ <= 8'H7e;
		32'H00210002: READ <= 8'H7e;
		32'H00210003: READ <= 8'H7f;
		32'H00210004: READ <= 8'H80;
		32'H00210005: READ <= 8'H80;
		32'H00210006: READ <= 8'H81;
		32'H00210007: READ <= 8'H82;
		32'H00210008: READ <= 8'H84;
		32'H00210009: READ <= 8'H86;
		32'H0021000a: READ <= 8'H88;
		32'H0021000b: READ <= 8'H8d;
		32'H0021000c: READ <= 8'H90;
		32'H0021000d: READ <= 8'H93;
		32'H0021000e: READ <= 8'H97;
		32'H0021000f: READ <= 8'H9b;
		32'H00210010: READ <= 8'H9e;
		32'H00210011: READ <= 8'Ha3;
		32'H00210012: READ <= 8'Hae;
		32'H00210013: READ <= 8'Hc9;
		32'H00210014: READ <= 8'Hcf;
		32'H00210015: READ <= 8'H99;
		32'H00210016: READ <= 8'H71;
		32'H00210017: READ <= 8'H68;
		32'H00210018: READ <= 8'H68;
		32'H00210019: READ <= 8'H65;
		32'H0021001a: READ <= 8'H64;
		32'H0021001b: READ <= 8'H68;
		32'H0021001c: READ <= 8'H5d;
		32'H0021001d: READ <= 8'H57;
		32'H0021001e: READ <= 8'H5e;
		32'H0021001f: READ <= 8'H64;
		32'H00210020: READ <= 8'H60;
		32'H00210021: READ <= 8'H33;
		32'H00210022: READ <= 8'H17;
		32'H00210023: READ <= 8'H1d;
		32'H00210024: READ <= 8'Hb;
		32'H00210025: READ <= 8'Ha;
		32'H00210026: READ <= 8'H4;
		32'H00210027: READ <= 8'H8;
		32'H00210028: READ <= 8'H49;
		32'H00210029: READ <= 8'H4d;
		32'H0021002a: READ <= 8'H52;
		32'H0021002b: READ <= 8'H59;
		32'H0021002c: READ <= 8'H4d;
		32'H0021002d: READ <= 8'H6d;
		32'H0021002e: READ <= 8'H6e;
		32'H0021002f: READ <= 8'H57;
		32'H00210030: READ <= 8'H63;
		32'H00210031: READ <= 8'H4b;
		32'H00210032: READ <= 8'H33;
		32'H00210033: READ <= 8'H2c;
		32'H00210034: READ <= 8'H4a;
		32'H00210035: READ <= 8'H5f;
		32'H00210036: READ <= 8'H1c;
		32'H00210037: READ <= 8'H3;
		32'H00210038: READ <= 8'H4;
		32'H00210039: READ <= 8'H22;
		32'H0021003a: READ <= 8'H74;
		32'H0021003b: READ <= 8'H75;
		32'H0021003c: READ <= 8'H91;
		32'H0021003d: READ <= 8'H97;
		32'H0021003e: READ <= 8'H9;
		32'H0021003f: READ <= 8'H6;
		32'H00210040: READ <= 8'H48;
		32'H00210041: READ <= 8'Ha0;
		32'H00210042: READ <= 8'H9b;
		32'H00210043: READ <= 8'Ha0;
		32'H00210044: READ <= 8'H9c;
		32'H00210045: READ <= 8'H98;
		32'H00210046: READ <= 8'H92;
		32'H00210047: READ <= 8'H8d;
		32'H00210048: READ <= 8'H90;
		32'H00210049: READ <= 8'H94;
		32'H0021004a: READ <= 8'H89;
		32'H0021004b: READ <= 8'H7d;
		32'H0021004c: READ <= 8'H59;
		32'H0021004d: READ <= 8'H71;
		32'H0021004e: READ <= 8'H82;
		32'H0021004f: READ <= 8'H89;
		32'H00210050: READ <= 8'H9c;
		32'H00210051: READ <= 8'H90;
		32'H00210052: READ <= 8'H9d;
		32'H00210053: READ <= 8'Hb1;
		32'H00210054: READ <= 8'Haf;
		32'H00210055: READ <= 8'H8a;
		32'H00210056: READ <= 8'H7c;
		32'H00210057: READ <= 8'H6f;
		32'H00210058: READ <= 8'H70;
		32'H00210059: READ <= 8'H79;
		32'H0021005a: READ <= 8'H85;
		32'H0021005b: READ <= 8'H85;
		32'H0021005c: READ <= 8'H85;
		32'H0021005d: READ <= 8'H85;
		32'H0021005e: READ <= 8'H86;
		32'H0021005f: READ <= 8'H87;
		32'H00210060: READ <= 8'H87;
		32'H00210061: READ <= 8'H87;
		32'H00210062: READ <= 8'H88;
		32'H00210063: READ <= 8'H88;
		
		32'H00220000: READ <= 8'H7c;
		32'H00220001: READ <= 8'H7d;
		32'H00220002: READ <= 8'H7d;
		32'H00220003: READ <= 8'H7e;
		32'H00220004: READ <= 8'H7e;
		32'H00220005: READ <= 8'H7f;
		32'H00220006: READ <= 8'H7f;
		32'H00220007: READ <= 8'H81;
		32'H00220008: READ <= 8'H81;
		32'H00220009: READ <= 8'H84;
		32'H0022000a: READ <= 8'H85;
		32'H0022000b: READ <= 8'H86;
		32'H0022000c: READ <= 8'H8b;
		32'H0022000d: READ <= 8'H90;
		32'H0022000e: READ <= 8'H93;
		32'H0022000f: READ <= 8'H96;
		32'H00220010: READ <= 8'H9a;
		32'H00220011: READ <= 8'Ha2;
		32'H00220012: READ <= 8'Hc2;
		32'H00220013: READ <= 8'Hdd;
		32'H00220014: READ <= 8'Hab;
		32'H00220015: READ <= 8'H84;
		32'H00220016: READ <= 8'H70;
		32'H00220017: READ <= 8'H50;
		32'H00220018: READ <= 8'H3b;
		32'H00220019: READ <= 8'H35;
		32'H0022001a: READ <= 8'H33;
		32'H0022001b: READ <= 8'H51;
		32'H0022001c: READ <= 8'H51;
		32'H0022001d: READ <= 8'H5f;
		32'H0022001e: READ <= 8'H4b;
		32'H0022001f: READ <= 8'H45;
		32'H00220020: READ <= 8'H47;
		32'H00220021: READ <= 8'H3b;
		32'H00220022: READ <= 8'H9;
		32'H00220023: READ <= 8'H13;
		32'H00220024: READ <= 8'H33;
		32'H00220025: READ <= 8'H1f;
		32'H00220026: READ <= 8'H10;
		32'H00220027: READ <= 8'H7;
		32'H00220028: READ <= 8'H15;
		32'H00220029: READ <= 8'H44;
		32'H0022002a: READ <= 8'H3b;
		32'H0022002b: READ <= 8'H50;
		32'H0022002c: READ <= 8'H58;
		32'H0022002d: READ <= 8'H3e;
		32'H0022002e: READ <= 8'H54;
		32'H0022002f: READ <= 8'H50;
		32'H00220030: READ <= 8'H71;
		32'H00220031: READ <= 8'H2e;
		32'H00220032: READ <= 8'H3e;
		32'H00220033: READ <= 8'H2c;
		32'H00220034: READ <= 8'H54;
		32'H00220035: READ <= 8'H4f;
		32'H00220036: READ <= 8'H17;
		32'H00220037: READ <= 8'H4;
		32'H00220038: READ <= 8'H3;
		32'H00220039: READ <= 8'H1f;
		32'H0022003a: READ <= 8'H6e;
		32'H0022003b: READ <= 8'H7b;
		32'H0022003c: READ <= 8'H93;
		32'H0022003d: READ <= 8'H92;
		32'H0022003e: READ <= 8'He;
		32'H0022003f: READ <= 8'Hd;
		32'H00220040: READ <= 8'H1c;
		32'H00220041: READ <= 8'H94;
		32'H00220042: READ <= 8'H98;
		32'H00220043: READ <= 8'H91;
		32'H00220044: READ <= 8'H93;
		32'H00220045: READ <= 8'H8e;
		32'H00220046: READ <= 8'H82;
		32'H00220047: READ <= 8'H8a;
		32'H00220048: READ <= 8'H91;
		32'H00220049: READ <= 8'H9b;
		32'H0022004a: READ <= 8'H86;
		32'H0022004b: READ <= 8'H7d;
		32'H0022004c: READ <= 8'H5e;
		32'H0022004d: READ <= 8'H68;
		32'H0022004e: READ <= 8'H84;
		32'H0022004f: READ <= 8'H80;
		32'H00220050: READ <= 8'H84;
		32'H00220051: READ <= 8'H85;
		32'H00220052: READ <= 8'H87;
		32'H00220053: READ <= 8'H8d;
		32'H00220054: READ <= 8'H94;
		32'H00220055: READ <= 8'H85;
		32'H00220056: READ <= 8'H92;
		32'H00220057: READ <= 8'H87;
		32'H00220058: READ <= 8'H84;
		32'H00220059: READ <= 8'H7a;
		32'H0022005a: READ <= 8'H7c;
		32'H0022005b: READ <= 8'H85;
		32'H0022005c: READ <= 8'H85;
		32'H0022005d: READ <= 8'H86;
		32'H0022005e: READ <= 8'H87;
		32'H0022005f: READ <= 8'H87;
		32'H00220060: READ <= 8'H87;
		32'H00220061: READ <= 8'H88;
		32'H00220062: READ <= 8'H88;
		32'H00220063: READ <= 8'H88;
		
		32'H00230000: READ <= 8'H7c;
		32'H00230001: READ <= 8'H7c;
		32'H00230002: READ <= 8'H7c;
		32'H00230003: READ <= 8'H7c;
		32'H00230004: READ <= 8'H7d;
		32'H00230005: READ <= 8'H7d;
		32'H00230006: READ <= 8'H7e;
		32'H00230007: READ <= 8'H80;
		32'H00230008: READ <= 8'H80;
		32'H00230009: READ <= 8'H81;
		32'H0023000a: READ <= 8'H83;
		32'H0023000b: READ <= 8'H83;
		32'H0023000c: READ <= 8'H86;
		32'H0023000d: READ <= 8'H8a;
		32'H0023000e: READ <= 8'H8e;
		32'H0023000f: READ <= 8'H92;
		32'H00230010: READ <= 8'H96;
		32'H00230011: READ <= 8'Ha2;
		32'H00230012: READ <= 8'Hc8;
		32'H00230013: READ <= 8'Hb6;
		32'H00230014: READ <= 8'H81;
		32'H00230015: READ <= 8'H6c;
		32'H00230016: READ <= 8'H6b;
		32'H00230017: READ <= 8'H3d;
		32'H00230018: READ <= 8'H20;
		32'H00230019: READ <= 8'H16;
		32'H0023001a: READ <= 8'H13;
		32'H0023001b: READ <= 8'H12;
		32'H0023001c: READ <= 8'H17;
		32'H0023001d: READ <= 8'H1a;
		32'H0023001e: READ <= 8'H1f;
		32'H0023001f: READ <= 8'H46;
		32'H00230020: READ <= 8'Hc;
		32'H00230021: READ <= 8'H11;
		32'H00230022: READ <= 8'H4;
		32'H00230023: READ <= 8'H2b;
		32'H00230024: READ <= 8'H37;
		32'H00230025: READ <= 8'H3a;
		32'H00230026: READ <= 8'H1e;
		32'H00230027: READ <= 8'H7;
		32'H00230028: READ <= 8'H7;
		32'H00230029: READ <= 8'H2e;
		32'H0023002a: READ <= 8'H64;
		32'H0023002b: READ <= 8'H32;
		32'H0023002c: READ <= 8'H60;
		32'H0023002d: READ <= 8'H5a;
		32'H0023002e: READ <= 8'H4b;
		32'H0023002f: READ <= 8'H57;
		32'H00230030: READ <= 8'H41;
		32'H00230031: READ <= 8'H4e;
		32'H00230032: READ <= 8'H3f;
		32'H00230033: READ <= 8'H20;
		32'H00230034: READ <= 8'H63;
		32'H00230035: READ <= 8'H4e;
		32'H00230036: READ <= 8'Hc;
		32'H00230037: READ <= 8'H4;
		32'H00230038: READ <= 8'Ha;
		32'H00230039: READ <= 8'H23;
		32'H0023003a: READ <= 8'H6c;
		32'H0023003b: READ <= 8'H77;
		32'H0023003c: READ <= 8'H8d;
		32'H0023003d: READ <= 8'H97;
		32'H0023003e: READ <= 8'H19;
		32'H0023003f: READ <= 8'H1a;
		32'H00230040: READ <= 8'Hf;
		32'H00230041: READ <= 8'H77;
		32'H00230042: READ <= 8'H8d;
		32'H00230043: READ <= 8'H90;
		32'H00230044: READ <= 8'H7f;
		32'H00230045: READ <= 8'H76;
		32'H00230046: READ <= 8'H7a;
		32'H00230047: READ <= 8'H92;
		32'H00230048: READ <= 8'H99;
		32'H00230049: READ <= 8'H9e;
		32'H0023004a: READ <= 8'H8c;
		32'H0023004b: READ <= 8'H80;
		32'H0023004c: READ <= 8'H70;
		32'H0023004d: READ <= 8'H63;
		32'H0023004e: READ <= 8'H7e;
		32'H0023004f: READ <= 8'H7f;
		32'H00230050: READ <= 8'H80;
		32'H00230051: READ <= 8'H81;
		32'H00230052: READ <= 8'H82;
		32'H00230053: READ <= 8'H82;
		32'H00230054: READ <= 8'H83;
		32'H00230055: READ <= 8'H85;
		32'H00230056: READ <= 8'H7a;
		32'H00230057: READ <= 8'H79;
		32'H00230058: READ <= 8'H8f;
		32'H00230059: READ <= 8'H89;
		32'H0023005a: READ <= 8'H88;
		32'H0023005b: READ <= 8'H85;
		32'H0023005c: READ <= 8'H86;
		32'H0023005d: READ <= 8'H86;
		32'H0023005e: READ <= 8'H87;
		32'H0023005f: READ <= 8'H87;
		32'H00230060: READ <= 8'H88;
		32'H00230061: READ <= 8'H87;
		32'H00230062: READ <= 8'H87;
		32'H00230063: READ <= 8'H88;
		
		32'H00240000: READ <= 8'H7b;
		32'H00240001: READ <= 8'H7a;
		32'H00240002: READ <= 8'H7b;
		32'H00240003: READ <= 8'H7b;
		32'H00240004: READ <= 8'H7b;
		32'H00240005: READ <= 8'H7c;
		32'H00240006: READ <= 8'H7d;
		32'H00240007: READ <= 8'H7e;
		32'H00240008: READ <= 8'H7f;
		32'H00240009: READ <= 8'H7f;
		32'H0024000a: READ <= 8'H81;
		32'H0024000b: READ <= 8'H81;
		32'H0024000c: READ <= 8'H82;
		32'H0024000d: READ <= 8'H86;
		32'H0024000e: READ <= 8'H89;
		32'H0024000f: READ <= 8'H8d;
		32'H00240010: READ <= 8'H91;
		32'H00240011: READ <= 8'Ha1;
		32'H00240012: READ <= 8'Hcc;
		32'H00240013: READ <= 8'Hac;
		32'H00240014: READ <= 8'H90;
		32'H00240015: READ <= 8'H56;
		32'H00240016: READ <= 8'H31;
		32'H00240017: READ <= 8'H28;
		32'H00240018: READ <= 8'H26;
		32'H00240019: READ <= 8'H2d;
		32'H0024001a: READ <= 8'H28;
		32'H0024001b: READ <= 8'H22;
		32'H0024001c: READ <= 8'H21;
		32'H0024001d: READ <= 8'H25;
		32'H0024001e: READ <= 8'H27;
		32'H0024001f: READ <= 8'H1d;
		32'H00240020: READ <= 8'H1c;
		32'H00240021: READ <= 8'H21;
		32'H00240022: READ <= 8'H18;
		32'H00240023: READ <= 8'H65;
		32'H00240024: READ <= 8'H6d;
		32'H00240025: READ <= 8'H30;
		32'H00240026: READ <= 8'H53;
		32'H00240027: READ <= 8'H2a;
		32'H00240028: READ <= 8'H8;
		32'H00240029: READ <= 8'H8;
		32'H0024002a: READ <= 8'H46;
		32'H0024002b: READ <= 8'H71;
		32'H0024002c: READ <= 8'H36;
		32'H0024002d: READ <= 8'H3e;
		32'H0024002e: READ <= 8'H48;
		32'H0024002f: READ <= 8'H49;
		32'H00240030: READ <= 8'H50;
		32'H00240031: READ <= 8'H31;
		32'H00240032: READ <= 8'H31;
		32'H00240033: READ <= 8'H2f;
		32'H00240034: READ <= 8'H53;
		32'H00240035: READ <= 8'H4b;
		32'H00240036: READ <= 8'Ha;
		32'H00240037: READ <= 8'H6;
		32'H00240038: READ <= 8'Ha;
		32'H00240039: READ <= 8'H22;
		32'H0024003a: READ <= 8'H5d;
		32'H0024003b: READ <= 8'H7e;
		32'H0024003c: READ <= 8'H8c;
		32'H0024003d: READ <= 8'H9e;
		32'H0024003e: READ <= 8'H1d;
		32'H0024003f: READ <= 8'H2a;
		32'H00240040: READ <= 8'H11;
		32'H00240041: READ <= 8'H5f;
		32'H00240042: READ <= 8'H7e;
		32'H00240043: READ <= 8'H6d;
		32'H00240044: READ <= 8'H6e;
		32'H00240045: READ <= 8'H76;
		32'H00240046: READ <= 8'H8a;
		32'H00240047: READ <= 8'H93;
		32'H00240048: READ <= 8'H96;
		32'H00240049: READ <= 8'H95;
		32'H0024004a: READ <= 8'H95;
		32'H0024004b: READ <= 8'H92;
		32'H0024004c: READ <= 8'H71;
		32'H0024004d: READ <= 8'H7e;
		32'H0024004e: READ <= 8'H85;
		32'H0024004f: READ <= 8'H7e;
		32'H00240050: READ <= 8'H7f;
		32'H00240051: READ <= 8'H7f;
		32'H00240052: READ <= 8'H80;
		32'H00240053: READ <= 8'H81;
		32'H00240054: READ <= 8'H81;
		32'H00240055: READ <= 8'H82;
		32'H00240056: READ <= 8'H86;
		32'H00240057: READ <= 8'H71;
		32'H00240058: READ <= 8'H8b;
		32'H00240059: READ <= 8'H91;
		32'H0024005a: READ <= 8'H85;
		32'H0024005b: READ <= 8'H83;
		32'H0024005c: READ <= 8'H86;
		32'H0024005d: READ <= 8'H86;
		32'H0024005e: READ <= 8'H87;
		32'H0024005f: READ <= 8'H87;
		32'H00240060: READ <= 8'H87;
		32'H00240061: READ <= 8'H87;
		32'H00240062: READ <= 8'H87;
		32'H00240063: READ <= 8'H88;
		
		32'H00250000: READ <= 8'H79;
		32'H00250001: READ <= 8'H79;
		32'H00250002: READ <= 8'H79;
		32'H00250003: READ <= 8'H79;
		32'H00250004: READ <= 8'H7a;
		32'H00250005: READ <= 8'H7b;
		32'H00250006: READ <= 8'H7c;
		32'H00250007: READ <= 8'H7d;
		32'H00250008: READ <= 8'H7e;
		32'H00250009: READ <= 8'H7e;
		32'H0025000a: READ <= 8'H7f;
		32'H0025000b: READ <= 8'H80;
		32'H0025000c: READ <= 8'H80;
		32'H0025000d: READ <= 8'H83;
		32'H0025000e: READ <= 8'H85;
		32'H0025000f: READ <= 8'H88;
		32'H00250010: READ <= 8'H90;
		32'H00250011: READ <= 8'Hb1;
		32'H00250012: READ <= 8'Hd1;
		32'H00250013: READ <= 8'Hb2;
		32'H00250014: READ <= 8'H89;
		32'H00250015: READ <= 8'H71;
		32'H00250016: READ <= 8'H4b;
		32'H00250017: READ <= 8'H27;
		32'H00250018: READ <= 8'H16;
		32'H00250019: READ <= 8'H13;
		32'H0025001a: READ <= 8'H14;
		32'H0025001b: READ <= 8'H1c;
		32'H0025001c: READ <= 8'H28;
		32'H0025001d: READ <= 8'H30;
		32'H0025001e: READ <= 8'H49;
		32'H0025001f: READ <= 8'H5c;
		32'H00250020: READ <= 8'H69;
		32'H00250021: READ <= 8'H63;
		32'H00250022: READ <= 8'H2b;
		32'H00250023: READ <= 8'H6f;
		32'H00250024: READ <= 8'H5e;
		32'H00250025: READ <= 8'H29;
		32'H00250026: READ <= 8'H4c;
		32'H00250027: READ <= 8'H71;
		32'H00250028: READ <= 8'H3c;
		32'H00250029: READ <= 8'H11;
		32'H0025002a: READ <= 8'H15;
		32'H0025002b: READ <= 8'H5e;
		32'H0025002c: READ <= 8'H61;
		32'H0025002d: READ <= 8'H55;
		32'H0025002e: READ <= 8'H56;
		32'H0025002f: READ <= 8'H55;
		32'H00250030: READ <= 8'H42;
		32'H00250031: READ <= 8'H32;
		32'H00250032: READ <= 8'H30;
		32'H00250033: READ <= 8'H40;
		32'H00250034: READ <= 8'H4e;
		32'H00250035: READ <= 8'H41;
		32'H00250036: READ <= 8'Hc;
		32'H00250037: READ <= 8'H5;
		32'H00250038: READ <= 8'H2;
		32'H00250039: READ <= 8'H1d;
		32'H0025003a: READ <= 8'H4a;
		32'H0025003b: READ <= 8'H80;
		32'H0025003c: READ <= 8'H80;
		32'H0025003d: READ <= 8'H9d;
		32'H0025003e: READ <= 8'H4d;
		32'H0025003f: READ <= 8'H4d;
		32'H00250040: READ <= 8'H1d;
		32'H00250041: READ <= 8'H59;
		32'H00250042: READ <= 8'H65;
		32'H00250043: READ <= 8'H70;
		32'H00250044: READ <= 8'H80;
		32'H00250045: READ <= 8'H80;
		32'H00250046: READ <= 8'H83;
		32'H00250047: READ <= 8'H94;
		32'H00250048: READ <= 8'H96;
		32'H00250049: READ <= 8'H99;
		32'H0025004a: READ <= 8'H9d;
		32'H0025004b: READ <= 8'H89;
		32'H0025004c: READ <= 8'H85;
		32'H0025004d: READ <= 8'H82;
		32'H0025004e: READ <= 8'H8a;
		32'H0025004f: READ <= 8'H7f;
		32'H00250050: READ <= 8'H7e;
		32'H00250051: READ <= 8'H7e;
		32'H00250052: READ <= 8'H7f;
		32'H00250053: READ <= 8'H80;
		32'H00250054: READ <= 8'H81;
		32'H00250055: READ <= 8'H81;
		32'H00250056: READ <= 8'H82;
		32'H00250057: READ <= 8'H85;
		32'H00250058: READ <= 8'H90;
		32'H00250059: READ <= 8'Ha2;
		32'H0025005a: READ <= 8'H97;
		32'H0025005b: READ <= 8'H86;
		32'H0025005c: READ <= 8'H85;
		32'H0025005d: READ <= 8'H86;
		32'H0025005e: READ <= 8'H87;
		32'H0025005f: READ <= 8'H86;
		32'H00250060: READ <= 8'H87;
		32'H00250061: READ <= 8'H87;
		32'H00250062: READ <= 8'H88;
		32'H00250063: READ <= 8'H88;
		
		32'H00260000: READ <= 8'H78;
		32'H00260001: READ <= 8'H78;
		32'H00260002: READ <= 8'H77;
		32'H00260003: READ <= 8'H78;
		32'H00260004: READ <= 8'H79;
		32'H00260005: READ <= 8'H79;
		32'H00260006: READ <= 8'H7b;
		32'H00260007: READ <= 8'H7c;
		32'H00260008: READ <= 8'H7c;
		32'H00260009: READ <= 8'H7d;
		32'H0026000a: READ <= 8'H7d;
		32'H0026000b: READ <= 8'H7d;
		32'H0026000c: READ <= 8'H7f;
		32'H0026000d: READ <= 8'H80;
		32'H0026000e: READ <= 8'H82;
		32'H0026000f: READ <= 8'H84;
		32'H00260010: READ <= 8'H89;
		32'H00260011: READ <= 8'Ha2;
		32'H00260012: READ <= 8'Hca;
		32'H00260013: READ <= 8'Hb2;
		32'H00260014: READ <= 8'H91;
		32'H00260015: READ <= 8'H74;
		32'H00260016: READ <= 8'H73;
		32'H00260017: READ <= 8'H54;
		32'H00260018: READ <= 8'H4d;
		32'H00260019: READ <= 8'H43;
		32'H0026001a: READ <= 8'H44;
		32'H0026001b: READ <= 8'H4d;
		32'H0026001c: READ <= 8'H61;
		32'H0026001d: READ <= 8'H66;
		32'H0026001e: READ <= 8'H75;
		32'H0026001f: READ <= 8'H73;
		32'H00260020: READ <= 8'H79;
		32'H00260021: READ <= 8'H64;
		32'H00260022: READ <= 8'H2e;
		32'H00260023: READ <= 8'H5e;
		32'H00260024: READ <= 8'H66;
		32'H00260025: READ <= 8'H57;
		32'H00260026: READ <= 8'H47;
		32'H00260027: READ <= 8'H6c;
		32'H00260028: READ <= 8'H7b;
		32'H00260029: READ <= 8'H55;
		32'H0026002a: READ <= 8'H13;
		32'H0026002b: READ <= 8'H19;
		32'H0026002c: READ <= 8'H59;
		32'H0026002d: READ <= 8'H4f;
		32'H0026002e: READ <= 8'H42;
		32'H0026002f: READ <= 8'H4a;
		32'H00260030: READ <= 8'H46;
		32'H00260031: READ <= 8'H43;
		32'H00260032: READ <= 8'H30;
		32'H00260033: READ <= 8'H53;
		32'H00260034: READ <= 8'H5d;
		32'H00260035: READ <= 8'H24;
		32'H00260036: READ <= 8'H19;
		32'H00260037: READ <= 8'H20;
		32'H00260038: READ <= 8'H7;
		32'H00260039: READ <= 8'H23;
		32'H0026003a: READ <= 8'H43;
		32'H0026003b: READ <= 8'H7a;
		32'H0026003c: READ <= 8'H77;
		32'H0026003d: READ <= 8'H91;
		32'H0026003e: READ <= 8'H6f;
		32'H0026003f: READ <= 8'H68;
		32'H00260040: READ <= 8'H2c;
		32'H00260041: READ <= 8'H6f;
		32'H00260042: READ <= 8'H5e;
		32'H00260043: READ <= 8'H7a;
		32'H00260044: READ <= 8'H8b;
		32'H00260045: READ <= 8'H86;
		32'H00260046: READ <= 8'H8b;
		32'H00260047: READ <= 8'H8b;
		32'H00260048: READ <= 8'H8a;
		32'H00260049: READ <= 8'H9a;
		32'H0026004a: READ <= 8'Ha4;
		32'H0026004b: READ <= 8'H8f;
		32'H0026004c: READ <= 8'H81;
		32'H0026004d: READ <= 8'H98;
		32'H0026004e: READ <= 8'H8f;
		32'H0026004f: READ <= 8'H7e;
		32'H00260050: READ <= 8'H7d;
		32'H00260051: READ <= 8'H7e;
		32'H00260052: READ <= 8'H7e;
		32'H00260053: READ <= 8'H7f;
		32'H00260054: READ <= 8'H80;
		32'H00260055: READ <= 8'H81;
		32'H00260056: READ <= 8'H82;
		32'H00260057: READ <= 8'H82;
		32'H00260058: READ <= 8'H8d;
		32'H00260059: READ <= 8'H9a;
		32'H0026005a: READ <= 8'Ha6;
		32'H0026005b: READ <= 8'H99;
		32'H0026005c: READ <= 8'H8a;
		32'H0026005d: READ <= 8'H86;
		32'H0026005e: READ <= 8'H86;
		32'H0026005f: READ <= 8'H87;
		32'H00260060: READ <= 8'H87;
		32'H00260061: READ <= 8'H87;
		32'H00260062: READ <= 8'H88;
		32'H00260063: READ <= 8'H88;
		
		32'H00270000: READ <= 8'H77;
		32'H00270001: READ <= 8'H77;
		32'H00270002: READ <= 8'H76;
		32'H00270003: READ <= 8'H77;
		32'H00270004: READ <= 8'H77;
		32'H00270005: READ <= 8'H79;
		32'H00270006: READ <= 8'H79;
		32'H00270007: READ <= 8'H7a;
		32'H00270008: READ <= 8'H7b;
		32'H00270009: READ <= 8'H7b;
		32'H0027000a: READ <= 8'H7b;
		32'H0027000b: READ <= 8'H7d;
		32'H0027000c: READ <= 8'H7d;
		32'H0027000d: READ <= 8'H7e;
		32'H0027000e: READ <= 8'H7f;
		32'H0027000f: READ <= 8'H81;
		32'H00270010: READ <= 8'H89;
		32'H00270011: READ <= 8'Haf;
		32'H00270012: READ <= 8'Hcf;
		32'H00270013: READ <= 8'Hb6;
		32'H00270014: READ <= 8'H7c;
		32'H00270015: READ <= 8'H86;
		32'H00270016: READ <= 8'H6a;
		32'H00270017: READ <= 8'H6b;
		32'H00270018: READ <= 8'H59;
		32'H00270019: READ <= 8'H4e;
		32'H0027001a: READ <= 8'H4d;
		32'H0027001b: READ <= 8'H51;
		32'H0027001c: READ <= 8'H62;
		32'H0027001d: READ <= 8'H76;
		32'H0027001e: READ <= 8'H70;
		32'H0027001f: READ <= 8'H71;
		32'H00270020: READ <= 8'H7d;
		32'H00270021: READ <= 8'H72;
		32'H00270022: READ <= 8'H37;
		32'H00270023: READ <= 8'H64;
		32'H00270024: READ <= 8'H6b;
		32'H00270025: READ <= 8'H6a;
		32'H00270026: READ <= 8'H35;
		32'H00270027: READ <= 8'H4a;
		32'H00270028: READ <= 8'H77;
		32'H00270029: READ <= 8'H77;
		32'H0027002a: READ <= 8'H4c;
		32'H0027002b: READ <= 8'H15;
		32'H0027002c: READ <= 8'H15;
		32'H0027002d: READ <= 8'H49;
		32'H0027002e: READ <= 8'H6c;
		32'H0027002f: READ <= 8'H3a;
		32'H00270030: READ <= 8'H35;
		32'H00270031: READ <= 8'H4b;
		32'H00270032: READ <= 8'H2e;
		32'H00270033: READ <= 8'H46;
		32'H00270034: READ <= 8'H6b;
		32'H00270035: READ <= 8'H8;
		32'H00270036: READ <= 8'H51;
		32'H00270037: READ <= 8'H94;
		32'H00270038: READ <= 8'H48;
		32'H00270039: READ <= 8'H33;
		32'H0027003a: READ <= 8'H36;
		32'H0027003b: READ <= 8'H70;
		32'H0027003c: READ <= 8'H70;
		32'H0027003d: READ <= 8'H92;
		32'H0027003e: READ <= 8'H72;
		32'H0027003f: READ <= 8'H6d;
		32'H00270040: READ <= 8'H33;
		32'H00270041: READ <= 8'H5d;
		32'H00270042: READ <= 8'H46;
		32'H00270043: READ <= 8'H6a;
		32'H00270044: READ <= 8'H8e;
		32'H00270045: READ <= 8'H7f;
		32'H00270046: READ <= 8'H81;
		32'H00270047: READ <= 8'H83;
		32'H00270048: READ <= 8'H8e;
		32'H00270049: READ <= 8'H92;
		32'H0027004a: READ <= 8'H99;
		32'H0027004b: READ <= 8'H94;
		32'H0027004c: READ <= 8'H88;
		32'H0027004d: READ <= 8'Ha5;
		32'H0027004e: READ <= 8'H97;
		32'H0027004f: READ <= 8'H7f;
		32'H00270050: READ <= 8'H7d;
		32'H00270051: READ <= 8'H7d;
		32'H00270052: READ <= 8'H7d;
		32'H00270053: READ <= 8'H7f;
		32'H00270054: READ <= 8'H7f;
		32'H00270055: READ <= 8'H80;
		32'H00270056: READ <= 8'H82;
		32'H00270057: READ <= 8'H82;
		32'H00270058: READ <= 8'H84;
		32'H00270059: READ <= 8'H92;
		32'H0027005a: READ <= 8'Ha1;
		32'H0027005b: READ <= 8'Ha8;
		32'H0027005c: READ <= 8'Ha0;
		32'H0027005d: READ <= 8'H8d;
		32'H0027005e: READ <= 8'H86;
		32'H0027005f: READ <= 8'H88;
		32'H00270060: READ <= 8'H87;
		32'H00270061: READ <= 8'H87;
		32'H00270062: READ <= 8'H88;
		32'H00270063: READ <= 8'H88;
		
		32'H00280000: READ <= 8'H76;
		32'H00280001: READ <= 8'H76;
		32'H00280002: READ <= 8'H75;
		32'H00280003: READ <= 8'H76;
		32'H00280004: READ <= 8'H76;
		32'H00280005: READ <= 8'H77;
		32'H00280006: READ <= 8'H77;
		32'H00280007: READ <= 8'H78;
		32'H00280008: READ <= 8'H79;
		32'H00280009: READ <= 8'H7a;
		32'H0028000a: READ <= 8'H7a;
		32'H0028000b: READ <= 8'H7b;
		32'H0028000c: READ <= 8'H7c;
		32'H0028000d: READ <= 8'H7c;
		32'H0028000e: READ <= 8'H7c;
		32'H0028000f: READ <= 8'H7f;
		32'H00280010: READ <= 8'H85;
		32'H00280011: READ <= 8'Ha9;
		32'H00280012: READ <= 8'Hc8;
		32'H00280013: READ <= 8'Hb0;
		32'H00280014: READ <= 8'H8c;
		32'H00280015: READ <= 8'H75;
		32'H00280016: READ <= 8'H69;
		32'H00280017: READ <= 8'H6e;
		32'H00280018: READ <= 8'H48;
		32'H00280019: READ <= 8'H4b;
		32'H0028001a: READ <= 8'H4c;
		32'H0028001b: READ <= 8'H5c;
		32'H0028001c: READ <= 8'H5a;
		32'H0028001d: READ <= 8'H6d;
		32'H0028001e: READ <= 8'H60;
		32'H0028001f: READ <= 8'H57;
		32'H00280020: READ <= 8'H60;
		32'H00280021: READ <= 8'H64;
		32'H00280022: READ <= 8'H3e;
		32'H00280023: READ <= 8'H61;
		32'H00280024: READ <= 8'H65;
		32'H00280025: READ <= 8'H6f;
		32'H00280026: READ <= 8'H48;
		32'H00280027: READ <= 8'H24;
		32'H00280028: READ <= 8'H60;
		32'H00280029: READ <= 8'H69;
		32'H0028002a: READ <= 8'H65;
		32'H0028002b: READ <= 8'H53;
		32'H0028002c: READ <= 8'H2a;
		32'H0028002d: READ <= 8'H1a;
		32'H0028002e: READ <= 8'H42;
		32'H0028002f: READ <= 8'H1c;
		32'H00280030: READ <= 8'H18;
		32'H00280031: READ <= 8'H34;
		32'H00280032: READ <= 8'H2a;
		32'H00280033: READ <= 8'H37;
		32'H00280034: READ <= 8'H5b;
		32'H00280035: READ <= 8'H3;
		32'H00280036: READ <= 8'H95;
		32'H00280037: READ <= 8'Hb7;
		32'H00280038: READ <= 8'Ha3;
		32'H00280039: READ <= 8'H6f;
		32'H0028003a: READ <= 8'H41;
		32'H0028003b: READ <= 8'H65;
		32'H0028003c: READ <= 8'H70;
		32'H0028003d: READ <= 8'H95;
		32'H0028003e: READ <= 8'H5d;
		32'H0028003f: READ <= 8'H5f;
		32'H00280040: READ <= 8'H46;
		32'H00280041: READ <= 8'H61;
		32'H00280042: READ <= 8'H5b;
		32'H00280043: READ <= 8'H5c;
		32'H00280044: READ <= 8'H7c;
		32'H00280045: READ <= 8'H81;
		32'H00280046: READ <= 8'H82;
		32'H00280047: READ <= 8'H89;
		32'H00280048: READ <= 8'H8d;
		32'H00280049: READ <= 8'H95;
		32'H0028004a: READ <= 8'H96;
		32'H0028004b: READ <= 8'H93;
		32'H0028004c: READ <= 8'H93;
		32'H0028004d: READ <= 8'Ha2;
		32'H0028004e: READ <= 8'H94;
		32'H0028004f: READ <= 8'H7f;
		32'H00280050: READ <= 8'H7c;
		32'H00280051: READ <= 8'H7c;
		32'H00280052: READ <= 8'H7d;
		32'H00280053: READ <= 8'H7e;
		32'H00280054: READ <= 8'H7f;
		32'H00280055: READ <= 8'H80;
		32'H00280056: READ <= 8'H81;
		32'H00280057: READ <= 8'H82;
		32'H00280058: READ <= 8'H82;
		32'H00280059: READ <= 8'H88;
		32'H0028005a: READ <= 8'H9f;
		32'H0028005b: READ <= 8'Ha5;
		32'H0028005c: READ <= 8'Haf;
		32'H0028005d: READ <= 8'Ha9;
		32'H0028005e: READ <= 8'H93;
		32'H0028005f: READ <= 8'H88;
		32'H00280060: READ <= 8'H88;
		32'H00280061: READ <= 8'H88;
		32'H00280062: READ <= 8'H88;
		32'H00280063: READ <= 8'H88;
		
		32'H00290000: READ <= 8'H75;
		32'H00290001: READ <= 8'H75;
		32'H00290002: READ <= 8'H74;
		32'H00290003: READ <= 8'H75;
		32'H00290004: READ <= 8'H75;
		32'H00290005: READ <= 8'H76;
		32'H00290006: READ <= 8'H77;
		32'H00290007: READ <= 8'H76;
		32'H00290008: READ <= 8'H77;
		32'H00290009: READ <= 8'H78;
		32'H0029000a: READ <= 8'H79;
		32'H0029000b: READ <= 8'H79;
		32'H0029000c: READ <= 8'H7a;
		32'H0029000d: READ <= 8'H7a;
		32'H0029000e: READ <= 8'H7c;
		32'H0029000f: READ <= 8'H7c;
		32'H00290010: READ <= 8'H81;
		32'H00290011: READ <= 8'H9a;
		32'H00290012: READ <= 8'Hbc;
		32'H00290013: READ <= 8'Ha8;
		32'H00290014: READ <= 8'H8c;
		32'H00290015: READ <= 8'H7d;
		32'H00290016: READ <= 8'H68;
		32'H00290017: READ <= 8'H62;
		32'H00290018: READ <= 8'H58;
		32'H00290019: READ <= 8'H53;
		32'H0029001a: READ <= 8'H4e;
		32'H0029001b: READ <= 8'H63;
		32'H0029001c: READ <= 8'H5d;
		32'H0029001d: READ <= 8'H5e;
		32'H0029001e: READ <= 8'H68;
		32'H0029001f: READ <= 8'H5e;
		32'H00290020: READ <= 8'H74;
		32'H00290021: READ <= 8'H69;
		32'H00290022: READ <= 8'H55;
		32'H00290023: READ <= 8'H42;
		32'H00290024: READ <= 8'H5c;
		32'H00290025: READ <= 8'H61;
		32'H00290026: READ <= 8'H60;
		32'H00290027: READ <= 8'H1e;
		32'H00290028: READ <= 8'H3a;
		32'H00290029: READ <= 8'H59;
		32'H0029002a: READ <= 8'H53;
		32'H0029002b: READ <= 8'H62;
		32'H0029002c: READ <= 8'H5e;
		32'H0029002d: READ <= 8'H1b;
		32'H0029002e: READ <= 8'He;
		32'H0029002f: READ <= 8'H3;
		32'H00290030: READ <= 8'H6;
		32'H00290031: READ <= 8'H23;
		32'H00290032: READ <= 8'H21;
		32'H00290033: READ <= 8'H1e;
		32'H00290034: READ <= 8'H2c;
		32'H00290035: READ <= 8'H51;
		32'H00290036: READ <= 8'Hdb;
		32'H00290037: READ <= 8'Ha9;
		32'H00290038: READ <= 8'H8a;
		32'H00290039: READ <= 8'H8a;
		32'H0029003a: READ <= 8'H44;
		32'H0029003b: READ <= 8'H60;
		32'H0029003c: READ <= 8'H6c;
		32'H0029003d: READ <= 8'H90;
		32'H0029003e: READ <= 8'H49;
		32'H0029003f: READ <= 8'H4c;
		32'H00290040: READ <= 8'H49;
		32'H00290041: READ <= 8'H69;
		32'H00290042: READ <= 8'H71;
		32'H00290043: READ <= 8'H66;
		32'H00290044: READ <= 8'H77;
		32'H00290045: READ <= 8'H76;
		32'H00290046: READ <= 8'H7b;
		32'H00290047: READ <= 8'H81;
		32'H00290048: READ <= 8'H85;
		32'H00290049: READ <= 8'H91;
		32'H0029004a: READ <= 8'H9b;
		32'H0029004b: READ <= 8'H99;
		32'H0029004c: READ <= 8'Ha1;
		32'H0029004d: READ <= 8'Ha8;
		32'H0029004e: READ <= 8'H97;
		32'H0029004f: READ <= 8'H7e;
		32'H00290050: READ <= 8'H7c;
		32'H00290051: READ <= 8'H7c;
		32'H00290052: READ <= 8'H7d;
		32'H00290053: READ <= 8'H7e;
		32'H00290054: READ <= 8'H7f;
		32'H00290055: READ <= 8'H7f;
		32'H00290056: READ <= 8'H80;
		32'H00290057: READ <= 8'H82;
		32'H00290058: READ <= 8'H82;
		32'H00290059: READ <= 8'H83;
		32'H0029005a: READ <= 8'H8f;
		32'H0029005b: READ <= 8'H9c;
		32'H0029005c: READ <= 8'H96;
		32'H0029005d: READ <= 8'Ha3;
		32'H0029005e: READ <= 8'H95;
		32'H0029005f: READ <= 8'H88;
		32'H00290060: READ <= 8'H88;
		32'H00290061: READ <= 8'H89;
		32'H00290062: READ <= 8'H88;
		32'H00290063: READ <= 8'H89;
		
		32'H002a0000: READ <= 8'H74;
		32'H002a0001: READ <= 8'H74;
		32'H002a0002: READ <= 8'H74;
		32'H002a0003: READ <= 8'H75;
		32'H002a0004: READ <= 8'H74;
		32'H002a0005: READ <= 8'H76;
		32'H002a0006: READ <= 8'H76;
		32'H002a0007: READ <= 8'H75;
		32'H002a0008: READ <= 8'H76;
		32'H002a0009: READ <= 8'H76;
		32'H002a000a: READ <= 8'H77;
		32'H002a000b: READ <= 8'H78;
		32'H002a000c: READ <= 8'H78;
		32'H002a000d: READ <= 8'H79;
		32'H002a000e: READ <= 8'H7a;
		32'H002a000f: READ <= 8'H7b;
		32'H002a0010: READ <= 8'H7d;
		32'H002a0011: READ <= 8'H95;
		32'H002a0012: READ <= 8'Hbc;
		32'H002a0013: READ <= 8'Hb0;
		32'H002a0014: READ <= 8'H89;
		32'H002a0015: READ <= 8'H6f;
		32'H002a0016: READ <= 8'H7a;
		32'H002a0017: READ <= 8'H6f;
		32'H002a0018: READ <= 8'H4e;
		32'H002a0019: READ <= 8'H48;
		32'H002a001a: READ <= 8'H3f;
		32'H002a001b: READ <= 8'H52;
		32'H002a001c: READ <= 8'H56;
		32'H002a001d: READ <= 8'H4d;
		32'H002a001e: READ <= 8'H4d;
		32'H002a001f: READ <= 8'H57;
		32'H002a0020: READ <= 8'H60;
		32'H002a0021: READ <= 8'H4f;
		32'H002a0022: READ <= 8'H3c;
		32'H002a0023: READ <= 8'H32;
		32'H002a0024: READ <= 8'H55;
		32'H002a0025: READ <= 8'H56;
		32'H002a0026: READ <= 8'H64;
		32'H002a0027: READ <= 8'H1a;
		32'H002a0028: READ <= 8'H1d;
		32'H002a0029: READ <= 8'H4e;
		32'H002a002a: READ <= 8'H59;
		32'H002a002b: READ <= 8'H47;
		32'H002a002c: READ <= 8'H42;
		32'H002a002d: READ <= 8'H23;
		32'H002a002e: READ <= 8'H18;
		32'H002a002f: READ <= 8'H8;
		32'H002a0030: READ <= 8'H11;
		32'H002a0031: READ <= 8'H31;
		32'H002a0032: READ <= 8'H33;
		32'H002a0033: READ <= 8'H9;
		32'H002a0034: READ <= 8'H1e;
		32'H002a0035: READ <= 8'Hcd;
		32'H002a0036: READ <= 8'Hfc;
		32'H002a0037: READ <= 8'Ha4;
		32'H002a0038: READ <= 8'H66;
		32'H002a0039: READ <= 8'H76;
		32'H002a003a: READ <= 8'H3a;
		32'H002a003b: READ <= 8'H5b;
		32'H002a003c: READ <= 8'H69;
		32'H002a003d: READ <= 8'H7e;
		32'H002a003e: READ <= 8'H30;
		32'H002a003f: READ <= 8'H3d;
		32'H002a0040: READ <= 8'H47;
		32'H002a0041: READ <= 8'H5d;
		32'H002a0042: READ <= 8'H68;
		32'H002a0043: READ <= 8'H6b;
		32'H002a0044: READ <= 8'H6c;
		32'H002a0045: READ <= 8'H69;
		32'H002a0046: READ <= 8'H6f;
		32'H002a0047: READ <= 8'H6c;
		32'H002a0048: READ <= 8'H88;
		32'H002a0049: READ <= 8'H8e;
		32'H002a004a: READ <= 8'H9d;
		32'H002a004b: READ <= 8'Ha9;
		32'H002a004c: READ <= 8'Ha4;
		32'H002a004d: READ <= 8'Ha8;
		32'H002a004e: READ <= 8'H9e;
		32'H002a004f: READ <= 8'H80;
		32'H002a0050: READ <= 8'H7b;
		32'H002a0051: READ <= 8'H7c;
		32'H002a0052: READ <= 8'H7c;
		32'H002a0053: READ <= 8'H7d;
		32'H002a0054: READ <= 8'H7e;
		32'H002a0055: READ <= 8'H7f;
		32'H002a0056: READ <= 8'H81;
		32'H002a0057: READ <= 8'H82;
		32'H002a0058: READ <= 8'H82;
		32'H002a0059: READ <= 8'H83;
		32'H002a005a: READ <= 8'H83;
		32'H002a005b: READ <= 8'H8a;
		32'H002a005c: READ <= 8'H86;
		32'H002a005d: READ <= 8'H8a;
		32'H002a005e: READ <= 8'H89;
		32'H002a005f: READ <= 8'H88;
		32'H002a0060: READ <= 8'H88;
		32'H002a0061: READ <= 8'H88;
		32'H002a0062: READ <= 8'H89;
		32'H002a0063: READ <= 8'H89;
		
		32'H002b0000: READ <= 8'H74;
		32'H002b0001: READ <= 8'H73;
		32'H002b0002: READ <= 8'H73;
		32'H002b0003: READ <= 8'H74;
		32'H002b0004: READ <= 8'H74;
		32'H002b0005: READ <= 8'H75;
		32'H002b0006: READ <= 8'H75;
		32'H002b0007: READ <= 8'H75;
		32'H002b0008: READ <= 8'H74;
		32'H002b0009: READ <= 8'H75;
		32'H002b000a: READ <= 8'H75;
		32'H002b000b: READ <= 8'H76;
		32'H002b000c: READ <= 8'H76;
		32'H002b000d: READ <= 8'H77;
		32'H002b000e: READ <= 8'H78;
		32'H002b000f: READ <= 8'H79;
		32'H002b0010: READ <= 8'H81;
		32'H002b0011: READ <= 8'H9e;
		32'H002b0012: READ <= 8'Hc3;
		32'H002b0013: READ <= 8'Hbd;
		32'H002b0014: READ <= 8'H89;
		32'H002b0015: READ <= 8'H51;
		32'H002b0016: READ <= 8'H79;
		32'H002b0017: READ <= 8'H6f;
		32'H002b0018: READ <= 8'H53;
		32'H002b0019: READ <= 8'H46;
		32'H002b001a: READ <= 8'H35;
		32'H002b001b: READ <= 8'H36;
		32'H002b001c: READ <= 8'H30;
		32'H002b001d: READ <= 8'H2e;
		32'H002b001e: READ <= 8'H30;
		32'H002b001f: READ <= 8'H34;
		32'H002b0020: READ <= 8'H2e;
		32'H002b0021: READ <= 8'H38;
		32'H002b0022: READ <= 8'H35;
		32'H002b0023: READ <= 8'H2b;
		32'H002b0024: READ <= 8'H4a;
		32'H002b0025: READ <= 8'H56;
		32'H002b0026: READ <= 8'H50;
		32'H002b0027: READ <= 8'H2a;
		32'H002b0028: READ <= 8'H10;
		32'H002b0029: READ <= 8'H37;
		32'H002b002a: READ <= 8'H52;
		32'H002b002b: READ <= 8'H36;
		32'H002b002c: READ <= 8'H1e;
		32'H002b002d: READ <= 8'H17;
		32'H002b002e: READ <= 8'H1a;
		32'H002b002f: READ <= 8'Hf;
		32'H002b0030: READ <= 8'H40;
		32'H002b0031: READ <= 8'H50;
		32'H002b0032: READ <= 8'H36;
		32'H002b0033: READ <= 8'H1;
		32'H002b0034: READ <= 8'H2a;
		32'H002b0035: READ <= 8'He6;
		32'H002b0036: READ <= 8'Hf7;
		32'H002b0037: READ <= 8'Hb5;
		32'H002b0038: READ <= 8'H5b;
		32'H002b0039: READ <= 8'H75;
		32'H002b003a: READ <= 8'H36;
		32'H002b003b: READ <= 8'H51;
		32'H002b003c: READ <= 8'H6c;
		32'H002b003d: READ <= 8'H76;
		32'H002b003e: READ <= 8'H1c;
		32'H002b003f: READ <= 8'H36;
		32'H002b0040: READ <= 8'H4a;
		32'H002b0041: READ <= 8'H5c;
		32'H002b0042: READ <= 8'H68;
		32'H002b0043: READ <= 8'H67;
		32'H002b0044: READ <= 8'H72;
		32'H002b0045: READ <= 8'H6e;
		32'H002b0046: READ <= 8'H69;
		32'H002b0047: READ <= 8'H69;
		32'H002b0048: READ <= 8'H84;
		32'H002b0049: READ <= 8'H90;
		32'H002b004a: READ <= 8'H98;
		32'H002b004b: READ <= 8'H97;
		32'H002b004c: READ <= 8'Ha7;
		32'H002b004d: READ <= 8'Hb3;
		32'H002b004e: READ <= 8'H9c;
		32'H002b004f: READ <= 8'H7f;
		32'H002b0050: READ <= 8'H7c;
		32'H002b0051: READ <= 8'H7b;
		32'H002b0052: READ <= 8'H7d;
		32'H002b0053: READ <= 8'H7d;
		32'H002b0054: READ <= 8'H7e;
		32'H002b0055: READ <= 8'H7f;
		32'H002b0056: READ <= 8'H81;
		32'H002b0057: READ <= 8'H81;
		32'H002b0058: READ <= 8'H82;
		32'H002b0059: READ <= 8'H83;
		32'H002b005a: READ <= 8'H84;
		32'H002b005b: READ <= 8'H85;
		32'H002b005c: READ <= 8'H86;
		32'H002b005d: READ <= 8'H87;
		32'H002b005e: READ <= 8'H88;
		32'H002b005f: READ <= 8'H88;
		32'H002b0060: READ <= 8'H88;
		32'H002b0061: READ <= 8'H89;
		32'H002b0062: READ <= 8'H89;
		32'H002b0063: READ <= 8'H88;
		
		32'H002c0000: READ <= 8'H73;
		32'H002c0001: READ <= 8'H73;
		32'H002c0002: READ <= 8'H73;
		32'H002c0003: READ <= 8'H73;
		32'H002c0004: READ <= 8'H73;
		32'H002c0005: READ <= 8'H74;
		32'H002c0006: READ <= 8'H75;
		32'H002c0007: READ <= 8'H75;
		32'H002c0008: READ <= 8'H74;
		32'H002c0009: READ <= 8'H74;
		32'H002c000a: READ <= 8'H74;
		32'H002c000b: READ <= 8'H75;
		32'H002c000c: READ <= 8'H75;
		32'H002c000d: READ <= 8'H76;
		32'H002c000e: READ <= 8'H77;
		32'H002c000f: READ <= 8'H78;
		32'H002c0010: READ <= 8'H7c;
		32'H002c0011: READ <= 8'H8e;
		32'H002c0012: READ <= 8'Hcb;
		32'H002c0013: READ <= 8'Hc7;
		32'H002c0014: READ <= 8'H91;
		32'H002c0015: READ <= 8'H57;
		32'H002c0016: READ <= 8'H6a;
		32'H002c0017: READ <= 8'H63;
		32'H002c0018: READ <= 8'H61;
		32'H002c0019: READ <= 8'H37;
		32'H002c001a: READ <= 8'H3f;
		32'H002c001b: READ <= 8'H3d;
		32'H002c001c: READ <= 8'H39;
		32'H002c001d: READ <= 8'H34;
		32'H002c001e: READ <= 8'H34;
		32'H002c001f: READ <= 8'H41;
		32'H002c0020: READ <= 8'H44;
		32'H002c0021: READ <= 8'H34;
		32'H002c0022: READ <= 8'H20;
		32'H002c0023: READ <= 8'H16;
		32'H002c0024: READ <= 8'H48;
		32'H002c0025: READ <= 8'H54;
		32'H002c0026: READ <= 8'H44;
		32'H002c0027: READ <= 8'H47;
		32'H002c0028: READ <= 8'H8;
		32'H002c0029: READ <= 8'H26;
		32'H002c002a: READ <= 8'H42;
		32'H002c002b: READ <= 8'H2d;
		32'H002c002c: READ <= 8'H18;
		32'H002c002d: READ <= 8'He;
		32'H002c002e: READ <= 8'H19;
		32'H002c002f: READ <= 8'H42;
		32'H002c0030: READ <= 8'H48;
		32'H002c0031: READ <= 8'H71;
		32'H002c0032: READ <= 8'H21;
		32'H002c0033: READ <= 8'H23;
		32'H002c0034: READ <= 8'H9e;
		32'H002c0035: READ <= 8'Hda;
		32'H002c0036: READ <= 8'He6;
		32'H002c0037: READ <= 8'Hca;
		32'H002c0038: READ <= 8'H6c;
		32'H002c0039: READ <= 8'H5f;
		32'H002c003a: READ <= 8'H2a;
		32'H002c003b: READ <= 8'H4f;
		32'H002c003c: READ <= 8'H6b;
		32'H002c003d: READ <= 8'H7c;
		32'H002c003e: READ <= 8'H24;
		32'H002c003f: READ <= 8'H2f;
		32'H002c0040: READ <= 8'H41;
		32'H002c0041: READ <= 8'H5b;
		32'H002c0042: READ <= 8'H62;
		32'H002c0043: READ <= 8'H65;
		32'H002c0044: READ <= 8'H65;
		32'H002c0045: READ <= 8'H62;
		32'H002c0046: READ <= 8'H75;
		32'H002c0047: READ <= 8'H71;
		32'H002c0048: READ <= 8'H90;
		32'H002c0049: READ <= 8'H94;
		32'H002c004a: READ <= 8'H9d;
		32'H002c004b: READ <= 8'Ha6;
		32'H002c004c: READ <= 8'Ha2;
		32'H002c004d: READ <= 8'Hb0;
		32'H002c004e: READ <= 8'H96;
		32'H002c004f: READ <= 8'H7e;
		32'H002c0050: READ <= 8'H7b;
		32'H002c0051: READ <= 8'H7b;
		32'H002c0052: READ <= 8'H7d;
		32'H002c0053: READ <= 8'H7e;
		32'H002c0054: READ <= 8'H7e;
		32'H002c0055: READ <= 8'H7f;
		32'H002c0056: READ <= 8'H81;
		32'H002c0057: READ <= 8'H81;
		32'H002c0058: READ <= 8'H82;
		32'H002c0059: READ <= 8'H83;
		32'H002c005a: READ <= 8'H84;
		32'H002c005b: READ <= 8'H85;
		32'H002c005c: READ <= 8'H86;
		32'H002c005d: READ <= 8'H86;
		32'H002c005e: READ <= 8'H88;
		32'H002c005f: READ <= 8'H88;
		32'H002c0060: READ <= 8'H88;
		32'H002c0061: READ <= 8'H89;
		32'H002c0062: READ <= 8'H89;
		32'H002c0063: READ <= 8'H89;
		
		32'H002d0000: READ <= 8'H73;
		32'H002d0001: READ <= 8'H72;
		32'H002d0002: READ <= 8'H72;
		32'H002d0003: READ <= 8'H73;
		32'H002d0004: READ <= 8'H73;
		32'H002d0005: READ <= 8'H74;
		32'H002d0006: READ <= 8'H75;
		32'H002d0007: READ <= 8'H74;
		32'H002d0008: READ <= 8'H74;
		32'H002d0009: READ <= 8'H74;
		32'H002d000a: READ <= 8'H74;
		32'H002d000b: READ <= 8'H74;
		32'H002d000c: READ <= 8'H74;
		32'H002d000d: READ <= 8'H75;
		32'H002d000e: READ <= 8'H76;
		32'H002d000f: READ <= 8'H78;
		32'H002d0010: READ <= 8'H80;
		32'H002d0011: READ <= 8'H9e;
		32'H002d0012: READ <= 8'Hbd;
		32'H002d0013: READ <= 8'Hb8;
		32'H002d0014: READ <= 8'Hae;
		32'H002d0015: READ <= 8'H83;
		32'H002d0016: READ <= 8'H78;
		32'H002d0017: READ <= 8'H6b;
		32'H002d0018: READ <= 8'H57;
		32'H002d0019: READ <= 8'H4a;
		32'H002d001a: READ <= 8'H48;
		32'H002d001b: READ <= 8'H3a;
		32'H002d001c: READ <= 8'H30;
		32'H002d001d: READ <= 8'H24;
		32'H002d001e: READ <= 8'H1c;
		32'H002d001f: READ <= 8'H1a;
		32'H002d0020: READ <= 8'H26;
		32'H002d0021: READ <= 8'H2f;
		32'H002d0022: READ <= 8'H2d;
		32'H002d0023: READ <= 8'Hc;
		32'H002d0024: READ <= 8'H37;
		32'H002d0025: READ <= 8'H48;
		32'H002d0026: READ <= 8'H33;
		32'H002d0027: READ <= 8'H4c;
		32'H002d0028: READ <= 8'Hc;
		32'H002d0029: READ <= 8'H16;
		32'H002d002a: READ <= 8'H2e;
		32'H002d002b: READ <= 8'H34;
		32'H002d002c: READ <= 8'H1e;
		32'H002d002d: READ <= 8'H26;
		32'H002d002e: READ <= 8'H6f;
		32'H002d002f: READ <= 8'Ha1;
		32'H002d0030: READ <= 8'Ha0;
		32'H002d0031: READ <= 8'H8d;
		32'H002d0032: READ <= 8'H4d;
		32'H002d0033: READ <= 8'H68;
		32'H002d0034: READ <= 8'Ha5;
		32'H002d0035: READ <= 8'Hc9;
		32'H002d0036: READ <= 8'Hd1;
		32'H002d0037: READ <= 8'Hca;
		32'H002d0038: READ <= 8'H78;
		32'H002d0039: READ <= 8'H4f;
		32'H002d003a: READ <= 8'H18;
		32'H002d003b: READ <= 8'H46;
		32'H002d003c: READ <= 8'H6b;
		32'H002d003d: READ <= 8'H88;
		32'H002d003e: READ <= 8'H43;
		32'H002d003f: READ <= 8'H36;
		32'H002d0040: READ <= 8'H4c;
		32'H002d0041: READ <= 8'H59;
		32'H002d0042: READ <= 8'H5e;
		32'H002d0043: READ <= 8'H6f;
		32'H002d0044: READ <= 8'H62;
		32'H002d0045: READ <= 8'H6e;
		32'H002d0046: READ <= 8'H72;
		32'H002d0047: READ <= 8'H71;
		32'H002d0048: READ <= 8'H7f;
		32'H002d0049: READ <= 8'H8a;
		32'H002d004a: READ <= 8'H92;
		32'H002d004b: READ <= 8'H9a;
		32'H002d004c: READ <= 8'Hac;
		32'H002d004d: READ <= 8'Had;
		32'H002d004e: READ <= 8'H93;
		32'H002d004f: READ <= 8'H7d;
		32'H002d0050: READ <= 8'H7b;
		32'H002d0051: READ <= 8'H7b;
		32'H002d0052: READ <= 8'H7c;
		32'H002d0053: READ <= 8'H7d;
		32'H002d0054: READ <= 8'H7e;
		32'H002d0055: READ <= 8'H7f;
		32'H002d0056: READ <= 8'H81;
		32'H002d0057: READ <= 8'H82;
		32'H002d0058: READ <= 8'H82;
		32'H002d0059: READ <= 8'H83;
		32'H002d005a: READ <= 8'H84;
		32'H002d005b: READ <= 8'H85;
		32'H002d005c: READ <= 8'H86;
		32'H002d005d: READ <= 8'H86;
		32'H002d005e: READ <= 8'H88;
		32'H002d005f: READ <= 8'H89;
		32'H002d0060: READ <= 8'H89;
		32'H002d0061: READ <= 8'H89;
		32'H002d0062: READ <= 8'H89;
		32'H002d0063: READ <= 8'H89;
		
		32'H002e0000: READ <= 8'H72;
		32'H002e0001: READ <= 8'H72;
		32'H002e0002: READ <= 8'H71;
		32'H002e0003: READ <= 8'H72;
		32'H002e0004: READ <= 8'H72;
		32'H002e0005: READ <= 8'H73;
		32'H002e0006: READ <= 8'H74;
		32'H002e0007: READ <= 8'H74;
		32'H002e0008: READ <= 8'H73;
		32'H002e0009: READ <= 8'H73;
		32'H002e000a: READ <= 8'H73;
		32'H002e000b: READ <= 8'H74;
		32'H002e000c: READ <= 8'H74;
		32'H002e000d: READ <= 8'H74;
		32'H002e000e: READ <= 8'H76;
		32'H002e000f: READ <= 8'H77;
		32'H002e0010: READ <= 8'H7a;
		32'H002e0011: READ <= 8'H89;
		32'H002e0012: READ <= 8'H9f;
		32'H002e0013: READ <= 8'Ha0;
		32'H002e0014: READ <= 8'Hb1;
		32'H002e0015: READ <= 8'H90;
		32'H002e0016: READ <= 8'H86;
		32'H002e0017: READ <= 8'H6c;
		32'H002e0018: READ <= 8'H51;
		32'H002e0019: READ <= 8'H54;
		32'H002e001a: READ <= 8'H47;
		32'H002e001b: READ <= 8'H35;
		32'H002e001c: READ <= 8'H2c;
		32'H002e001d: READ <= 8'H22;
		32'H002e001e: READ <= 8'H1a;
		32'H002e001f: READ <= 8'H16;
		32'H002e0020: READ <= 8'H15;
		32'H002e0021: READ <= 8'H15;
		32'H002e0022: READ <= 8'H14;
		32'H002e0023: READ <= 8'Hb;
		32'H002e0024: READ <= 8'H27;
		32'H002e0025: READ <= 8'H43;
		32'H002e0026: READ <= 8'H1c;
		32'H002e0027: READ <= 8'H50;
		32'H002e0028: READ <= 8'He;
		32'H002e0029: READ <= 8'Hd;
		32'H002e002a: READ <= 8'H17;
		32'H002e002b: READ <= 8'H30;
		32'H002e002c: READ <= 8'H5f;
		32'H002e002d: READ <= 8'Hc3;
		32'H002e002e: READ <= 8'Hef;
		32'H002e002f: READ <= 8'Hf1;
		32'H002e0030: READ <= 8'Hda;
		32'H002e0031: READ <= 8'Hb7;
		32'H002e0032: READ <= 8'Haf;
		32'H002e0033: READ <= 8'H9a;
		32'H002e0034: READ <= 8'Ha1;
		32'H002e0035: READ <= 8'Hb3;
		32'H002e0036: READ <= 8'Hb4;
		32'H002e0037: READ <= 8'Hbe;
		32'H002e0038: READ <= 8'H82;
		32'H002e0039: READ <= 8'H59;
		32'H002e003a: READ <= 8'H2f;
		32'H002e003b: READ <= 8'H26;
		32'H002e003c: READ <= 8'H54;
		32'H002e003d: READ <= 8'H8f;
		32'H002e003e: READ <= 8'H61;
		32'H002e003f: READ <= 8'H5d;
		32'H002e0040: READ <= 8'H3c;
		32'H002e0041: READ <= 8'H56;
		32'H002e0042: READ <= 8'H6d;
		32'H002e0043: READ <= 8'H6c;
		32'H002e0044: READ <= 8'H7f;
		32'H002e0045: READ <= 8'H71;
		32'H002e0046: READ <= 8'H7e;
		32'H002e0047: READ <= 8'H85;
		32'H002e0048: READ <= 8'H8b;
		32'H002e0049: READ <= 8'H92;
		32'H002e004a: READ <= 8'H9c;
		32'H002e004b: READ <= 8'Ha1;
		32'H002e004c: READ <= 8'H9f;
		32'H002e004d: READ <= 8'Ha9;
		32'H002e004e: READ <= 8'H8c;
		32'H002e004f: READ <= 8'H7b;
		32'H002e0050: READ <= 8'H7a;
		32'H002e0051: READ <= 8'H7b;
		32'H002e0052: READ <= 8'H7c;
		32'H002e0053: READ <= 8'H7d;
		32'H002e0054: READ <= 8'H7d;
		32'H002e0055: READ <= 8'H7f;
		32'H002e0056: READ <= 8'H80;
		32'H002e0057: READ <= 8'H81;
		32'H002e0058: READ <= 8'H82;
		32'H002e0059: READ <= 8'H83;
		32'H002e005a: READ <= 8'H84;
		32'H002e005b: READ <= 8'H85;
		32'H002e005c: READ <= 8'H86;
		32'H002e005d: READ <= 8'H87;
		32'H002e005e: READ <= 8'H89;
		32'H002e005f: READ <= 8'H89;
		32'H002e0060: READ <= 8'H89;
		32'H002e0061: READ <= 8'H89;
		32'H002e0062: READ <= 8'H8a;
		32'H002e0063: READ <= 8'H8a;
		
		32'H002f0000: READ <= 8'H71;
		32'H002f0001: READ <= 8'H71;
		32'H002f0002: READ <= 8'H71;
		32'H002f0003: READ <= 8'H71;
		32'H002f0004: READ <= 8'H72;
		32'H002f0005: READ <= 8'H72;
		32'H002f0006: READ <= 8'H73;
		32'H002f0007: READ <= 8'H73;
		32'H002f0008: READ <= 8'H73;
		32'H002f0009: READ <= 8'H73;
		32'H002f000a: READ <= 8'H73;
		32'H002f000b: READ <= 8'H73;
		32'H002f000c: READ <= 8'H73;
		32'H002f000d: READ <= 8'H74;
		32'H002f000e: READ <= 8'H74;
		32'H002f000f: READ <= 8'H75;
		32'H002f0010: READ <= 8'H78;
		32'H002f0011: READ <= 8'H82;
		32'H002f0012: READ <= 8'H85;
		32'H002f0013: READ <= 8'Ha6;
		32'H002f0014: READ <= 8'Hb9;
		32'H002f0015: READ <= 8'Hc3;
		32'H002f0016: READ <= 8'Ha5;
		32'H002f0017: READ <= 8'H83;
		32'H002f0018: READ <= 8'H61;
		32'H002f0019: READ <= 8'H5b;
		32'H002f001a: READ <= 8'H45;
		32'H002f001b: READ <= 8'H2d;
		32'H002f001c: READ <= 8'H27;
		32'H002f001d: READ <= 8'H22;
		32'H002f001e: READ <= 8'H1d;
		32'H002f001f: READ <= 8'H1a;
		32'H002f0020: READ <= 8'H16;
		32'H002f0021: READ <= 8'He;
		32'H002f0022: READ <= 8'Ha;
		32'H002f0023: READ <= 8'H6;
		32'H002f0024: READ <= 8'H20;
		32'H002f0025: READ <= 8'H44;
		32'H002f0026: READ <= 8'H26;
		32'H002f0027: READ <= 8'H50;
		32'H002f0028: READ <= 8'H1e;
		32'H002f0029: READ <= 8'H15;
		32'H002f002a: READ <= 8'H26;
		32'H002f002b: READ <= 8'H3a;
		32'H002f002c: READ <= 8'Hbb;
		32'H002f002d: READ <= 8'Hea;
		32'H002f002e: READ <= 8'Hea;
		32'H002f002f: READ <= 8'He5;
		32'H002f0030: READ <= 8'He6;
		32'H002f0031: READ <= 8'He0;
		32'H002f0032: READ <= 8'Hd2;
		32'H002f0033: READ <= 8'Hc5;
		32'H002f0034: READ <= 8'Hb9;
		32'H002f0035: READ <= 8'Ha5;
		32'H002f0036: READ <= 8'Ha8;
		32'H002f0037: READ <= 8'Ha4;
		32'H002f0038: READ <= 8'H8e;
		32'H002f0039: READ <= 8'H7a;
		32'H002f003a: READ <= 8'H74;
		32'H002f003b: READ <= 8'H3a;
		32'H002f003c: READ <= 8'H34;
		32'H002f003d: READ <= 8'H7c;
		32'H002f003e: READ <= 8'H74;
		32'H002f003f: READ <= 8'H72;
		32'H002f0040: READ <= 8'H3a;
		32'H002f0041: READ <= 8'H5d;
		32'H002f0042: READ <= 8'H62;
		32'H002f0043: READ <= 8'H64;
		32'H002f0044: READ <= 8'H73;
		32'H002f0045: READ <= 8'H77;
		32'H002f0046: READ <= 8'H81;
		32'H002f0047: READ <= 8'H83;
		32'H002f0048: READ <= 8'H84;
		32'H002f0049: READ <= 8'H90;
		32'H002f004a: READ <= 8'H9a;
		32'H002f004b: READ <= 8'H9e;
		32'H002f004c: READ <= 8'Hb1;
		32'H002f004d: READ <= 8'H98;
		32'H002f004e: READ <= 8'H88;
		32'H002f004f: READ <= 8'H7b;
		32'H002f0050: READ <= 8'H7b;
		32'H002f0051: READ <= 8'H7b;
		32'H002f0052: READ <= 8'H7c;
		32'H002f0053: READ <= 8'H7d;
		32'H002f0054: READ <= 8'H7d;
		32'H002f0055: READ <= 8'H7f;
		32'H002f0056: READ <= 8'H81;
		32'H002f0057: READ <= 8'H81;
		32'H002f0058: READ <= 8'H82;
		32'H002f0059: READ <= 8'H83;
		32'H002f005a: READ <= 8'H84;
		32'H002f005b: READ <= 8'H85;
		32'H002f005c: READ <= 8'H86;
		32'H002f005d: READ <= 8'H87;
		32'H002f005e: READ <= 8'H88;
		32'H002f005f: READ <= 8'H88;
		32'H002f0060: READ <= 8'H89;
		32'H002f0061: READ <= 8'H89;
		32'H002f0062: READ <= 8'H89;
		32'H002f0063: READ <= 8'H8a;
		
		32'H00300000: READ <= 8'H71;
		32'H00300001: READ <= 8'H71;
		32'H00300002: READ <= 8'H71;
		32'H00300003: READ <= 8'H70;
		32'H00300004: READ <= 8'H71;
		32'H00300005: READ <= 8'H71;
		32'H00300006: READ <= 8'H72;
		32'H00300007: READ <= 8'H73;
		32'H00300008: READ <= 8'H73;
		32'H00300009: READ <= 8'H72;
		32'H0030000a: READ <= 8'H72;
		32'H0030000b: READ <= 8'H72;
		32'H0030000c: READ <= 8'H72;
		32'H0030000d: READ <= 8'H73;
		32'H0030000e: READ <= 8'H73;
		32'H0030000f: READ <= 8'H74;
		32'H00300010: READ <= 8'H75;
		32'H00300011: READ <= 8'H77;
		32'H00300012: READ <= 8'H82;
		32'H00300013: READ <= 8'H90;
		32'H00300014: READ <= 8'Had;
		32'H00300015: READ <= 8'Hbe;
		32'H00300016: READ <= 8'Hbc;
		32'H00300017: READ <= 8'H99;
		32'H00300018: READ <= 8'H65;
		32'H00300019: READ <= 8'H60;
		32'H0030001a: READ <= 8'H51;
		32'H0030001b: READ <= 8'H22;
		32'H0030001c: READ <= 8'H20;
		32'H0030001d: READ <= 8'H1f;
		32'H0030001e: READ <= 8'H1e;
		32'H0030001f: READ <= 8'H1c;
		32'H00300020: READ <= 8'H18;
		32'H00300021: READ <= 8'Hf;
		32'H00300022: READ <= 8'H9;
		32'H00300023: READ <= 8'H7;
		32'H00300024: READ <= 8'He;
		32'H00300025: READ <= 8'H48;
		32'H00300026: READ <= 8'H2e;
		32'H00300027: READ <= 8'H4c;
		32'H00300028: READ <= 8'H44;
		32'H00300029: READ <= 8'H21;
		32'H0030002a: READ <= 8'H33;
		32'H0030002b: READ <= 8'H8f;
		32'H0030002c: READ <= 8'He1;
		32'H0030002d: READ <= 8'He2;
		32'H0030002e: READ <= 8'Hdb;
		32'H0030002f: READ <= 8'Hd8;
		32'H00300030: READ <= 8'Hdf;
		32'H00300031: READ <= 8'He2;
		32'H00300032: READ <= 8'Hdd;
		32'H00300033: READ <= 8'Hdc;
		32'H00300034: READ <= 8'Hcc;
		32'H00300035: READ <= 8'Hb0;
		32'H00300036: READ <= 8'Ha1;
		32'H00300037: READ <= 8'Ha3;
		32'H00300038: READ <= 8'H9e;
		32'H00300039: READ <= 8'H86;
		32'H0030003a: READ <= 8'H8e;
		32'H0030003b: READ <= 8'H37;
		32'H0030003c: READ <= 8'H5a;
		32'H0030003d: READ <= 8'H87;
		32'H0030003e: READ <= 8'H8c;
		32'H0030003f: READ <= 8'H71;
		32'H00300040: READ <= 8'H34;
		32'H00300041: READ <= 8'H62;
		32'H00300042: READ <= 8'H64;
		32'H00300043: READ <= 8'H71;
		32'H00300044: READ <= 8'H66;
		32'H00300045: READ <= 8'H75;
		32'H00300046: READ <= 8'H80;
		32'H00300047: READ <= 8'H81;
		32'H00300048: READ <= 8'H85;
		32'H00300049: READ <= 8'H99;
		32'H0030004a: READ <= 8'H9d;
		32'H0030004b: READ <= 8'Hab;
		32'H0030004c: READ <= 8'Haa;
		32'H0030004d: READ <= 8'H90;
		32'H0030004e: READ <= 8'H81;
		32'H0030004f: READ <= 8'H7b;
		32'H00300050: READ <= 8'H7b;
		32'H00300051: READ <= 8'H7b;
		32'H00300052: READ <= 8'H7c;
		32'H00300053: READ <= 8'H7d;
		32'H00300054: READ <= 8'H7e;
		32'H00300055: READ <= 8'H7f;
		32'H00300056: READ <= 8'H80;
		32'H00300057: READ <= 8'H81;
		32'H00300058: READ <= 8'H82;
		32'H00300059: READ <= 8'H83;
		32'H0030005a: READ <= 8'H84;
		32'H0030005b: READ <= 8'H85;
		32'H0030005c: READ <= 8'H86;
		32'H0030005d: READ <= 8'H87;
		32'H0030005e: READ <= 8'H89;
		32'H0030005f: READ <= 8'H88;
		32'H00300060: READ <= 8'H89;
		32'H00300061: READ <= 8'H89;
		32'H00300062: READ <= 8'H8a;
		32'H00300063: READ <= 8'H8a;
		
		32'H00310000: READ <= 8'H70;
		32'H00310001: READ <= 8'H70;
		32'H00310002: READ <= 8'H70;
		32'H00310003: READ <= 8'H70;
		32'H00310004: READ <= 8'H70;
		32'H00310005: READ <= 8'H71;
		32'H00310006: READ <= 8'H71;
		32'H00310007: READ <= 8'H71;
		32'H00310008: READ <= 8'H72;
		32'H00310009: READ <= 8'H72;
		32'H0031000a: READ <= 8'H72;
		32'H0031000b: READ <= 8'H71;
		32'H0031000c: READ <= 8'H71;
		32'H0031000d: READ <= 8'H71;
		32'H0031000e: READ <= 8'H72;
		32'H0031000f: READ <= 8'H73;
		32'H00310010: READ <= 8'H74;
		32'H00310011: READ <= 8'H76;
		32'H00310012: READ <= 8'H79;
		32'H00310013: READ <= 8'H7f;
		32'H00310014: READ <= 8'H97;
		32'H00310015: READ <= 8'Had;
		32'H00310016: READ <= 8'Hb7;
		32'H00310017: READ <= 8'Hb7;
		32'H00310018: READ <= 8'H91;
		32'H00310019: READ <= 8'H69;
		32'H0031001a: READ <= 8'H66;
		32'H0031001b: READ <= 8'H3c;
		32'H0031001c: READ <= 8'H1e;
		32'H0031001d: READ <= 8'H1c;
		32'H0031001e: READ <= 8'H20;
		32'H0031001f: READ <= 8'H20;
		32'H00310020: READ <= 8'H19;
		32'H00310021: READ <= 8'He;
		32'H00310022: READ <= 8'H8;
		32'H00310023: READ <= 8'H6;
		32'H00310024: READ <= 8'Hb;
		32'H00310025: READ <= 8'H40;
		32'H00310026: READ <= 8'H34;
		32'H00310027: READ <= 8'H50;
		32'H00310028: READ <= 8'H75;
		32'H00310029: READ <= 8'H3c;
		32'H0031002a: READ <= 8'H51;
		32'H0031002b: READ <= 8'Hc6;
		32'H0031002c: READ <= 8'Hcd;
		32'H0031002d: READ <= 8'Hd6;
		32'H0031002e: READ <= 8'Hd8;
		32'H0031002f: READ <= 8'Hdb;
		32'H00310030: READ <= 8'Hde;
		32'H00310031: READ <= 8'Hdb;
		32'H00310032: READ <= 8'Hd8;
		32'H00310033: READ <= 8'Hd6;
		32'H00310034: READ <= 8'Hc6;
		32'H00310035: READ <= 8'Hb3;
		32'H00310036: READ <= 8'Ha8;
		32'H00310037: READ <= 8'H9e;
		32'H00310038: READ <= 8'H9a;
		32'H00310039: READ <= 8'H8b;
		32'H0031003a: READ <= 8'H9a;
		32'H0031003b: READ <= 8'H45;
		32'H0031003c: READ <= 8'H65;
		32'H0031003d: READ <= 8'H9b;
		32'H0031003e: READ <= 8'H89;
		32'H0031003f: READ <= 8'H8c;
		32'H00310040: READ <= 8'H35;
		32'H00310041: READ <= 8'H4f;
		32'H00310042: READ <= 8'H59;
		32'H00310043: READ <= 8'H60;
		32'H00310044: READ <= 8'H63;
		32'H00310045: READ <= 8'H6f;
		32'H00310046: READ <= 8'H73;
		32'H00310047: READ <= 8'H83;
		32'H00310048: READ <= 8'H89;
		32'H00310049: READ <= 8'H99;
		32'H0031004a: READ <= 8'H9d;
		32'H0031004b: READ <= 8'Ha2;
		32'H0031004c: READ <= 8'H8e;
		32'H0031004d: READ <= 8'H84;
		32'H0031004e: READ <= 8'H7a;
		32'H0031004f: READ <= 8'H7b;
		32'H00310050: READ <= 8'H7b;
		32'H00310051: READ <= 8'H7c;
		32'H00310052: READ <= 8'H7d;
		32'H00310053: READ <= 8'H7d;
		32'H00310054: READ <= 8'H7e;
		32'H00310055: READ <= 8'H7f;
		32'H00310056: READ <= 8'H80;
		32'H00310057: READ <= 8'H81;
		32'H00310058: READ <= 8'H82;
		32'H00310059: READ <= 8'H82;
		32'H0031005a: READ <= 8'H84;
		32'H0031005b: READ <= 8'H84;
		32'H0031005c: READ <= 8'H86;
		32'H0031005d: READ <= 8'H87;
		32'H0031005e: READ <= 8'H88;
		32'H0031005f: READ <= 8'H88;
		32'H00310060: READ <= 8'H89;
		32'H00310061: READ <= 8'H89;
		32'H00310062: READ <= 8'H8a;
		32'H00310063: READ <= 8'H8a;
		
		32'H00320000: READ <= 8'H70;
		32'H00320001: READ <= 8'H70;
		32'H00320002: READ <= 8'H70;
		32'H00320003: READ <= 8'H70;
		32'H00320004: READ <= 8'H6f;
		32'H00320005: READ <= 8'H70;
		32'H00320006: READ <= 8'H70;
		32'H00320007: READ <= 8'H70;
		32'H00320008: READ <= 8'H71;
		32'H00320009: READ <= 8'H71;
		32'H0032000a: READ <= 8'H71;
		32'H0032000b: READ <= 8'H71;
		32'H0032000c: READ <= 8'H70;
		32'H0032000d: READ <= 8'H71;
		32'H0032000e: READ <= 8'H71;
		32'H0032000f: READ <= 8'H72;
		32'H00320010: READ <= 8'H73;
		32'H00320011: READ <= 8'H74;
		32'H00320012: READ <= 8'H77;
		32'H00320013: READ <= 8'H78;
		32'H00320014: READ <= 8'H87;
		32'H00320015: READ <= 8'H8e;
		32'H00320016: READ <= 8'H97;
		32'H00320017: READ <= 8'H96;
		32'H00320018: READ <= 8'Ha0;
		32'H00320019: READ <= 8'H8f;
		32'H0032001a: READ <= 8'H84;
		32'H0032001b: READ <= 8'H77;
		32'H0032001c: READ <= 8'H4a;
		32'H0032001d: READ <= 8'H2f;
		32'H0032001e: READ <= 8'H2a;
		32'H0032001f: READ <= 8'H27;
		32'H00320020: READ <= 8'H1d;
		32'H00320021: READ <= 8'H13;
		32'H00320022: READ <= 8'Hf;
		32'H00320023: READ <= 8'Hc;
		32'H00320024: READ <= 8'Hc;
		32'H00320025: READ <= 8'H2c;
		32'H00320026: READ <= 8'H29;
		32'H00320027: READ <= 8'H54;
		32'H00320028: READ <= 8'H4d;
		32'H00320029: READ <= 8'H61;
		32'H0032002a: READ <= 8'H85;
		32'H0032002b: READ <= 8'Hb2;
		32'H0032002c: READ <= 8'Hb9;
		32'H0032002d: READ <= 8'Hd4;
		32'H0032002e: READ <= 8'Hde;
		32'H0032002f: READ <= 8'He2;
		32'H00320030: READ <= 8'He7;
		32'H00320031: READ <= 8'He6;
		32'H00320032: READ <= 8'He0;
		32'H00320033: READ <= 8'Hd9;
		32'H00320034: READ <= 8'Hc9;
		32'H00320035: READ <= 8'Had;
		32'H00320036: READ <= 8'Hb2;
		32'H00320037: READ <= 8'H9b;
		32'H00320038: READ <= 8'H9e;
		32'H00320039: READ <= 8'H8f;
		32'H0032003a: READ <= 8'H9f;
		32'H0032003b: READ <= 8'H4f;
		32'H0032003c: READ <= 8'H52;
		32'H0032003d: READ <= 8'H9f;
		32'H0032003e: READ <= 8'H78;
		32'H0032003f: READ <= 8'Ha1;
		32'H00320040: READ <= 8'H37;
		32'H00320041: READ <= 8'H59;
		32'H00320042: READ <= 8'H5d;
		32'H00320043: READ <= 8'H6a;
		32'H00320044: READ <= 8'H65;
		32'H00320045: READ <= 8'H5d;
		32'H00320046: READ <= 8'H62;
		32'H00320047: READ <= 8'H67;
		32'H00320048: READ <= 8'H72;
		32'H00320049: READ <= 8'H84;
		32'H0032004a: READ <= 8'H8e;
		32'H0032004b: READ <= 8'H91;
		32'H0032004c: READ <= 8'H92;
		32'H0032004d: READ <= 8'H7c;
		32'H0032004e: READ <= 8'H7a;
		32'H0032004f: READ <= 8'H7a;
		32'H00320050: READ <= 8'H7a;
		32'H00320051: READ <= 8'H7b;
		32'H00320052: READ <= 8'H7c;
		32'H00320053: READ <= 8'H7e;
		32'H00320054: READ <= 8'H7e;
		32'H00320055: READ <= 8'H7f;
		32'H00320056: READ <= 8'H80;
		32'H00320057: READ <= 8'H81;
		32'H00320058: READ <= 8'H82;
		32'H00320059: READ <= 8'H83;
		32'H0032005a: READ <= 8'H83;
		32'H0032005b: READ <= 8'H85;
		32'H0032005c: READ <= 8'H86;
		32'H0032005d: READ <= 8'H87;
		32'H0032005e: READ <= 8'H88;
		32'H0032005f: READ <= 8'H89;
		32'H00320060: READ <= 8'H89;
		32'H00320061: READ <= 8'H8a;
		32'H00320062: READ <= 8'H8a;
		32'H00320063: READ <= 8'H89;
		
		32'H00330000: READ <= 8'H70;
		32'H00330001: READ <= 8'H6f;
		32'H00330002: READ <= 8'H6f;
		32'H00330003: READ <= 8'H6f;
		32'H00330004: READ <= 8'H70;
		32'H00330005: READ <= 8'H70;
		32'H00330006: READ <= 8'H70;
		32'H00330007: READ <= 8'H6f;
		32'H00330008: READ <= 8'H70;
		32'H00330009: READ <= 8'H70;
		32'H0033000a: READ <= 8'H70;
		32'H0033000b: READ <= 8'H71;
		32'H0033000c: READ <= 8'H6f;
		32'H0033000d: READ <= 8'H6f;
		32'H0033000e: READ <= 8'H70;
		32'H0033000f: READ <= 8'H71;
		32'H00330010: READ <= 8'H72;
		32'H00330011: READ <= 8'H74;
		32'H00330012: READ <= 8'H76;
		32'H00330013: READ <= 8'H78;
		32'H00330014: READ <= 8'H7b;
		32'H00330015: READ <= 8'H7d;
		32'H00330016: READ <= 8'H82;
		32'H00330017: READ <= 8'H87;
		32'H00330018: READ <= 8'H8c;
		32'H00330019: READ <= 8'H92;
		32'H0033001a: READ <= 8'H9e;
		32'H0033001b: READ <= 8'H8c;
		32'H0033001c: READ <= 8'H5d;
		32'H0033001d: READ <= 8'H4f;
		32'H0033001e: READ <= 8'H45;
		32'H0033001f: READ <= 8'H40;
		32'H00330020: READ <= 8'H31;
		32'H00330021: READ <= 8'H24;
		32'H00330022: READ <= 8'H19;
		32'H00330023: READ <= 8'Hf;
		32'H00330024: READ <= 8'H1f;
		32'H00330025: READ <= 8'H37;
		32'H00330026: READ <= 8'H34;
		32'H00330027: READ <= 8'H28;
		32'H00330028: READ <= 8'H29;
		32'H00330029: READ <= 8'H70;
		32'H0033002a: READ <= 8'H8d;
		32'H0033002b: READ <= 8'Ha2;
		32'H0033002c: READ <= 8'Hc1;
		32'H0033002d: READ <= 8'Hda;
		32'H0033002e: READ <= 8'He0;
		32'H0033002f: READ <= 8'He4;
		32'H00330030: READ <= 8'He9;
		32'H00330031: READ <= 8'Heb;
		32'H00330032: READ <= 8'He8;
		32'H00330033: READ <= 8'He1;
		32'H00330034: READ <= 8'Hd1;
		32'H00330035: READ <= 8'Hbc;
		32'H00330036: READ <= 8'Hbe;
		32'H00330037: READ <= 8'Hb2;
		32'H00330038: READ <= 8'H9a;
		32'H00330039: READ <= 8'H9d;
		32'H0033003a: READ <= 8'H9b;
		32'H0033003b: READ <= 8'H61;
		32'H0033003c: READ <= 8'H47;
		32'H0033003d: READ <= 8'Ha1;
		32'H0033003e: READ <= 8'H75;
		32'H0033003f: READ <= 8'H9b;
		32'H00330040: READ <= 8'H4a;
		32'H00330041: READ <= 8'H7a;
		32'H00330042: READ <= 8'H64;
		32'H00330043: READ <= 8'H64;
		32'H00330044: READ <= 8'H70;
		32'H00330045: READ <= 8'H73;
		32'H00330046: READ <= 8'H7f;
		32'H00330047: READ <= 8'H85;
		32'H00330048: READ <= 8'H91;
		32'H00330049: READ <= 8'Ha0;
		32'H0033004a: READ <= 8'Ha8;
		32'H0033004b: READ <= 8'Ha1;
		32'H0033004c: READ <= 8'H91;
		32'H0033004d: READ <= 8'H78;
		32'H0033004e: READ <= 8'H7a;
		32'H0033004f: READ <= 8'H7a;
		32'H00330050: READ <= 8'H7a;
		32'H00330051: READ <= 8'H7b;
		32'H00330052: READ <= 8'H7d;
		32'H00330053: READ <= 8'H7e;
		32'H00330054: READ <= 8'H7e;
		32'H00330055: READ <= 8'H7f;
		32'H00330056: READ <= 8'H80;
		32'H00330057: READ <= 8'H81;
		32'H00330058: READ <= 8'H81;
		32'H00330059: READ <= 8'H83;
		32'H0033005a: READ <= 8'H83;
		32'H0033005b: READ <= 8'H84;
		32'H0033005c: READ <= 8'H86;
		32'H0033005d: READ <= 8'H87;
		32'H0033005e: READ <= 8'H88;
		32'H0033005f: READ <= 8'H89;
		32'H00330060: READ <= 8'H89;
		32'H00330061: READ <= 8'H8a;
		32'H00330062: READ <= 8'H8a;
		32'H00330063: READ <= 8'H89;
		
		32'H00340000: READ <= 8'H70;
		32'H00340001: READ <= 8'H70;
		32'H00340002: READ <= 8'H6f;
		32'H00340003: READ <= 8'H6f;
		32'H00340004: READ <= 8'H6f;
		32'H00340005: READ <= 8'H6f;
		32'H00340006: READ <= 8'H6f;
		32'H00340007: READ <= 8'H6f;
		32'H00340008: READ <= 8'H6f;
		32'H00340009: READ <= 8'H70;
		32'H0034000a: READ <= 8'H6f;
		32'H0034000b: READ <= 8'H6f;
		32'H0034000c: READ <= 8'H6f;
		32'H0034000d: READ <= 8'H6f;
		32'H0034000e: READ <= 8'H6f;
		32'H0034000f: READ <= 8'H70;
		32'H00340010: READ <= 8'H71;
		32'H00340011: READ <= 8'H72;
		32'H00340012: READ <= 8'H73;
		32'H00340013: READ <= 8'H77;
		32'H00340014: READ <= 8'H78;
		32'H00340015: READ <= 8'H7a;
		32'H00340016: READ <= 8'H7e;
		32'H00340017: READ <= 8'H81;
		32'H00340018: READ <= 8'H86;
		32'H00340019: READ <= 8'H91;
		32'H0034001a: READ <= 8'H8b;
		32'H0034001b: READ <= 8'H57;
		32'H0034001c: READ <= 8'H55;
		32'H0034001d: READ <= 8'H57;
		32'H0034001e: READ <= 8'H31;
		32'H0034001f: READ <= 8'H1a;
		32'H00340020: READ <= 8'H1f;
		32'H00340021: READ <= 8'H12;
		32'H00340022: READ <= 8'Hf;
		32'H00340023: READ <= 8'H12;
		32'H00340024: READ <= 8'H16;
		32'H00340025: READ <= 8'H3f;
		32'H00340026: READ <= 8'H2d;
		32'H00340027: READ <= 8'H10;
		32'H00340028: READ <= 8'H56;
		32'H00340029: READ <= 8'H72;
		32'H0034002a: READ <= 8'H9c;
		32'H0034002b: READ <= 8'Hb7;
		32'H0034002c: READ <= 8'Hce;
		32'H0034002d: READ <= 8'Hde;
		32'H0034002e: READ <= 8'He2;
		32'H0034002f: READ <= 8'He5;
		32'H00340030: READ <= 8'He9;
		32'H00340031: READ <= 8'Heb;
		32'H00340032: READ <= 8'He9;
		32'H00340033: READ <= 8'He3;
		32'H00340034: READ <= 8'Hd1;
		32'H00340035: READ <= 8'Hc4;
		32'H00340036: READ <= 8'Hc9;
		32'H00340037: READ <= 8'Hb7;
		32'H00340038: READ <= 8'Ha6;
		32'H00340039: READ <= 8'H8c;
		32'H0034003a: READ <= 8'H90;
		32'H0034003b: READ <= 8'H71;
		32'H0034003c: READ <= 8'H33;
		32'H0034003d: READ <= 8'H9a;
		32'H0034003e: READ <= 8'H7c;
		32'H0034003f: READ <= 8'H98;
		32'H00340040: READ <= 8'H52;
		32'H00340041: READ <= 8'H78;
		32'H00340042: READ <= 8'H6c;
		32'H00340043: READ <= 8'H65;
		32'H00340044: READ <= 8'H77;
		32'H00340045: READ <= 8'H87;
		32'H00340046: READ <= 8'H83;
		32'H00340047: READ <= 8'H9a;
		32'H00340048: READ <= 8'Ha2;
		32'H00340049: READ <= 8'Ha8;
		32'H0034004a: READ <= 8'Hb1;
		32'H0034004b: READ <= 8'Ha5;
		32'H0034004c: READ <= 8'H7c;
		32'H0034004d: READ <= 8'H79;
		32'H0034004e: READ <= 8'H79;
		32'H0034004f: READ <= 8'H7a;
		32'H00340050: READ <= 8'H7b;
		32'H00340051: READ <= 8'H7b;
		32'H00340052: READ <= 8'H7c;
		32'H00340053: READ <= 8'H7d;
		32'H00340054: READ <= 8'H7e;
		32'H00340055: READ <= 8'H7f;
		32'H00340056: READ <= 8'H80;
		32'H00340057: READ <= 8'H80;
		32'H00340058: READ <= 8'H81;
		32'H00340059: READ <= 8'H82;
		32'H0034005a: READ <= 8'H84;
		32'H0034005b: READ <= 8'H85;
		32'H0034005c: READ <= 8'H86;
		32'H0034005d: READ <= 8'H87;
		32'H0034005e: READ <= 8'H87;
		32'H0034005f: READ <= 8'H89;
		32'H00340060: READ <= 8'H89;
		32'H00340061: READ <= 8'H89;
		32'H00340062: READ <= 8'H8a;
		32'H00340063: READ <= 8'H8a;
		
		32'H00350000: READ <= 8'H70;
		32'H00350001: READ <= 8'H70;
		32'H00350002: READ <= 8'H6f;
		32'H00350003: READ <= 8'H70;
		32'H00350004: READ <= 8'H6f;
		32'H00350005: READ <= 8'H6f;
		32'H00350006: READ <= 8'H6e;
		32'H00350007: READ <= 8'H6f;
		32'H00350008: READ <= 8'H6e;
		32'H00350009: READ <= 8'H6e;
		32'H0035000a: READ <= 8'H6e;
		32'H0035000b: READ <= 8'H6e;
		32'H0035000c: READ <= 8'H6e;
		32'H0035000d: READ <= 8'H6e;
		32'H0035000e: READ <= 8'H6e;
		32'H0035000f: READ <= 8'H6f;
		32'H00350010: READ <= 8'H70;
		32'H00350011: READ <= 8'H71;
		32'H00350012: READ <= 8'H73;
		32'H00350013: READ <= 8'H74;
		32'H00350014: READ <= 8'H76;
		32'H00350015: READ <= 8'H78;
		32'H00350016: READ <= 8'H7b;
		32'H00350017: READ <= 8'H7d;
		32'H00350018: READ <= 8'H7f;
		32'H00350019: READ <= 8'H85;
		32'H0035001a: READ <= 8'H65;
		32'H0035001b: READ <= 8'H45;
		32'H0035001c: READ <= 8'H52;
		32'H0035001d: READ <= 8'H32;
		32'H0035001e: READ <= 8'H5;
		32'H0035001f: READ <= 8'H9;
		32'H00350020: READ <= 8'Hf;
		32'H00350021: READ <= 8'Hf;
		32'H00350022: READ <= 8'He;
		32'H00350023: READ <= 8'Hd;
		32'H00350024: READ <= 8'H1f;
		32'H00350025: READ <= 8'H47;
		32'H00350026: READ <= 8'H3c;
		32'H00350027: READ <= 8'H58;
		32'H00350028: READ <= 8'H77;
		32'H00350029: READ <= 8'H7f;
		32'H0035002a: READ <= 8'Hb0;
		32'H0035002b: READ <= 8'Hc7;
		32'H0035002c: READ <= 8'Hd9;
		32'H0035002d: READ <= 8'He0;
		32'H0035002e: READ <= 8'He3;
		32'H0035002f: READ <= 8'He6;
		32'H00350030: READ <= 8'He9;
		32'H00350031: READ <= 8'Heb;
		32'H00350032: READ <= 8'He9;
		32'H00350033: READ <= 8'He2;
		32'H00350034: READ <= 8'Hd3;
		32'H00350035: READ <= 8'Hc9;
		32'H00350036: READ <= 8'Hca;
		32'H00350037: READ <= 8'Hb7;
		32'H00350038: READ <= 8'Ha7;
		32'H00350039: READ <= 8'H91;
		32'H0035003a: READ <= 8'H85;
		32'H0035003b: READ <= 8'H73;
		32'H0035003c: READ <= 8'H2d;
		32'H0035003d: READ <= 8'H93;
		32'H0035003e: READ <= 8'H7d;
		32'H0035003f: READ <= 8'H85;
		32'H00350040: READ <= 8'H57;
		32'H00350041: READ <= 8'H79;
		32'H00350042: READ <= 8'H77;
		32'H00350043: READ <= 8'H52;
		32'H00350044: READ <= 8'H65;
		32'H00350045: READ <= 8'H77;
		32'H00350046: READ <= 8'H93;
		32'H00350047: READ <= 8'H97;
		32'H00350048: READ <= 8'Ha0;
		32'H00350049: READ <= 8'Hb3;
		32'H0035004a: READ <= 8'Haa;
		32'H0035004b: READ <= 8'H96;
		32'H0035004c: READ <= 8'H78;
		32'H0035004d: READ <= 8'H79;
		32'H0035004e: READ <= 8'H79;
		32'H0035004f: READ <= 8'H7a;
		32'H00350050: READ <= 8'H7b;
		32'H00350051: READ <= 8'H7b;
		32'H00350052: READ <= 8'H7d;
		32'H00350053: READ <= 8'H7d;
		32'H00350054: READ <= 8'H7d;
		32'H00350055: READ <= 8'H7e;
		32'H00350056: READ <= 8'H80;
		32'H00350057: READ <= 8'H80;
		32'H00350058: READ <= 8'H81;
		32'H00350059: READ <= 8'H82;
		32'H0035005a: READ <= 8'H84;
		32'H0035005b: READ <= 8'H85;
		32'H0035005c: READ <= 8'H86;
		32'H0035005d: READ <= 8'H86;
		32'H0035005e: READ <= 8'H87;
		32'H0035005f: READ <= 8'H88;
		32'H00350060: READ <= 8'H89;
		32'H00350061: READ <= 8'H8a;
		32'H00350062: READ <= 8'H8a;
		32'H00350063: READ <= 8'H89;
		
		32'H00360000: READ <= 8'H70;
		32'H00360001: READ <= 8'H70;
		32'H00360002: READ <= 8'H6f;
		32'H00360003: READ <= 8'H6f;
		32'H00360004: READ <= 8'H6f;
		32'H00360005: READ <= 8'H6f;
		32'H00360006: READ <= 8'H6e;
		32'H00360007: READ <= 8'H6e;
		32'H00360008: READ <= 8'H6e;
		32'H00360009: READ <= 8'H6e;
		32'H0036000a: READ <= 8'H6d;
		32'H0036000b: READ <= 8'H6d;
		32'H0036000c: READ <= 8'H6d;
		32'H0036000d: READ <= 8'H6d;
		32'H0036000e: READ <= 8'H6e;
		32'H0036000f: READ <= 8'H6e;
		32'H00360010: READ <= 8'H6e;
		32'H00360011: READ <= 8'H70;
		32'H00360012: READ <= 8'H72;
		32'H00360013: READ <= 8'H74;
		32'H00360014: READ <= 8'H74;
		32'H00360015: READ <= 8'H77;
		32'H00360016: READ <= 8'H78;
		32'H00360017: READ <= 8'H7b;
		32'H00360018: READ <= 8'H7c;
		32'H00360019: READ <= 8'H81;
		32'H0036001a: READ <= 8'H5b;
		32'H0036001b: READ <= 8'H4c;
		32'H0036001c: READ <= 8'H5e;
		32'H0036001d: READ <= 8'Hc;
		32'H0036001e: READ <= 8'Hd;
		32'H0036001f: READ <= 8'H14;
		32'H00360020: READ <= 8'H16;
		32'H00360021: READ <= 8'H13;
		32'H00360022: READ <= 8'H1a;
		32'H00360023: READ <= 8'H1c;
		32'H00360024: READ <= 8'H5f;
		32'H00360025: READ <= 8'H45;
		32'H00360026: READ <= 8'H4d;
		32'H00360027: READ <= 8'H5e;
		32'H00360028: READ <= 8'H7e;
		32'H00360029: READ <= 8'Ha7;
		32'H0036002a: READ <= 8'Hc1;
		32'H0036002b: READ <= 8'Hd0;
		32'H0036002c: READ <= 8'Hdd;
		32'H0036002d: READ <= 8'He1;
		32'H0036002e: READ <= 8'He3;
		32'H0036002f: READ <= 8'He6;
		32'H00360030: READ <= 8'He8;
		32'H00360031: READ <= 8'He9;
		32'H00360032: READ <= 8'He7;
		32'H00360033: READ <= 8'He0;
		32'H00360034: READ <= 8'Hd5;
		32'H00360035: READ <= 8'Hd0;
		32'H00360036: READ <= 8'Hcd;
		32'H00360037: READ <= 8'Hc6;
		32'H00360038: READ <= 8'Hc3;
		32'H00360039: READ <= 8'Hb6;
		32'H0036003a: READ <= 8'H8b;
		32'H0036003b: READ <= 8'H75;
		32'H0036003c: READ <= 8'H16;
		32'H0036003d: READ <= 8'H94;
		32'H0036003e: READ <= 8'H82;
		32'H0036003f: READ <= 8'H76;
		32'H00360040: READ <= 8'H65;
		32'H00360041: READ <= 8'H7c;
		32'H00360042: READ <= 8'H64;
		32'H00360043: READ <= 8'H70;
		32'H00360044: READ <= 8'H78;
		32'H00360045: READ <= 8'H87;
		32'H00360046: READ <= 8'H8f;
		32'H00360047: READ <= 8'H99;
		32'H00360048: READ <= 8'Had;
		32'H00360049: READ <= 8'Hb0;
		32'H0036004a: READ <= 8'Ha9;
		32'H0036004b: READ <= 8'H83;
		32'H0036004c: READ <= 8'H78;
		32'H0036004d: READ <= 8'H79;
		32'H0036004e: READ <= 8'H79;
		32'H0036004f: READ <= 8'H7a;
		32'H00360050: READ <= 8'H7b;
		32'H00360051: READ <= 8'H7b;
		32'H00360052: READ <= 8'H7c;
		32'H00360053: READ <= 8'H7d;
		32'H00360054: READ <= 8'H7e;
		32'H00360055: READ <= 8'H7f;
		32'H00360056: READ <= 8'H80;
		32'H00360057: READ <= 8'H81;
		32'H00360058: READ <= 8'H81;
		32'H00360059: READ <= 8'H82;
		32'H0036005a: READ <= 8'H83;
		32'H0036005b: READ <= 8'H84;
		32'H0036005c: READ <= 8'H85;
		32'H0036005d: READ <= 8'H87;
		32'H0036005e: READ <= 8'H88;
		32'H0036005f: READ <= 8'H89;
		32'H00360060: READ <= 8'H89;
		32'H00360061: READ <= 8'H89;
		32'H00360062: READ <= 8'H89;
		32'H00360063: READ <= 8'H8a;
		
		32'H00370000: READ <= 8'H70;
		32'H00370001: READ <= 8'H70;
		32'H00370002: READ <= 8'H6f;
		32'H00370003: READ <= 8'H70;
		32'H00370004: READ <= 8'H70;
		32'H00370005: READ <= 8'H6f;
		32'H00370006: READ <= 8'H6e;
		32'H00370007: READ <= 8'H6d;
		32'H00370008: READ <= 8'H6e;
		32'H00370009: READ <= 8'H6d;
		32'H0037000a: READ <= 8'H6d;
		32'H0037000b: READ <= 8'H6d;
		32'H0037000c: READ <= 8'H6c;
		32'H0037000d: READ <= 8'H6c;
		32'H0037000e: READ <= 8'H6d;
		32'H0037000f: READ <= 8'H6d;
		32'H00370010: READ <= 8'H6d;
		32'H00370011: READ <= 8'H6f;
		32'H00370012: READ <= 8'H70;
		32'H00370013: READ <= 8'H72;
		32'H00370014: READ <= 8'H74;
		32'H00370015: READ <= 8'H74;
		32'H00370016: READ <= 8'H76;
		32'H00370017: READ <= 8'H78;
		32'H00370018: READ <= 8'H7a;
		32'H00370019: READ <= 8'H7b;
		32'H0037001a: READ <= 8'H82;
		32'H0037001b: READ <= 8'H8a;
		32'H0037001c: READ <= 8'H77;
		32'H0037001d: READ <= 8'H2f;
		32'H0037001e: READ <= 8'H30;
		32'H0037001f: READ <= 8'H24;
		32'H00370020: READ <= 8'H3f;
		32'H00370021: READ <= 8'H62;
		32'H00370022: READ <= 8'H7f;
		32'H00370023: READ <= 8'H86;
		32'H00370024: READ <= 8'H89;
		32'H00370025: READ <= 8'H47;
		32'H00370026: READ <= 8'H48;
		32'H00370027: READ <= 8'H4e;
		32'H00370028: READ <= 8'H7e;
		32'H00370029: READ <= 8'Hb6;
		32'H0037002a: READ <= 8'Hc9;
		32'H0037002b: READ <= 8'Hd5;
		32'H0037002c: READ <= 8'Hde;
		32'H0037002d: READ <= 8'He1;
		32'H0037002e: READ <= 8'He2;
		32'H0037002f: READ <= 8'He4;
		32'H00370030: READ <= 8'He6;
		32'H00370031: READ <= 8'He7;
		32'H00370032: READ <= 8'He5;
		32'H00370033: READ <= 8'Hde;
		32'H00370034: READ <= 8'Hd8;
		32'H00370035: READ <= 8'Hd4;
		32'H00370036: READ <= 8'Hd4;
		32'H00370037: READ <= 8'Hd3;
		32'H00370038: READ <= 8'Hd3;
		32'H00370039: READ <= 8'Hd4;
		32'H0037003a: READ <= 8'H9e;
		32'H0037003b: READ <= 8'H71;
		32'H0037003c: READ <= 8'H17;
		32'H0037003d: READ <= 8'H7e;
		32'H0037003e: READ <= 8'H87;
		32'H0037003f: READ <= 8'H6c;
		32'H00370040: READ <= 8'H6e;
		32'H00370041: READ <= 8'H73;
		32'H00370042: READ <= 8'H6c;
		32'H00370043: READ <= 8'H71;
		32'H00370044: READ <= 8'H7d;
		32'H00370045: READ <= 8'H8a;
		32'H00370046: READ <= 8'H98;
		32'H00370047: READ <= 8'H9b;
		32'H00370048: READ <= 8'Hb1;
		32'H00370049: READ <= 8'Haf;
		32'H0037004a: READ <= 8'H96;
		32'H0037004b: READ <= 8'H7c;
		32'H0037004c: READ <= 8'H78;
		32'H0037004d: READ <= 8'H78;
		32'H0037004e: READ <= 8'H7a;
		32'H0037004f: READ <= 8'H7a;
		32'H00370050: READ <= 8'H7a;
		32'H00370051: READ <= 8'H7b;
		32'H00370052: READ <= 8'H7c;
		32'H00370053: READ <= 8'H7d;
		32'H00370054: READ <= 8'H7e;
		32'H00370055: READ <= 8'H7e;
		32'H00370056: READ <= 8'H80;
		32'H00370057: READ <= 8'H81;
		32'H00370058: READ <= 8'H82;
		32'H00370059: READ <= 8'H82;
		32'H0037005a: READ <= 8'H84;
		32'H0037005b: READ <= 8'H84;
		32'H0037005c: READ <= 8'H86;
		32'H0037005d: READ <= 8'H87;
		32'H0037005e: READ <= 8'H88;
		32'H0037005f: READ <= 8'H89;
		32'H00370060: READ <= 8'H88;
		32'H00370061: READ <= 8'H89;
		32'H00370062: READ <= 8'H8a;
		32'H00370063: READ <= 8'H8a;
		
		32'H00380000: READ <= 8'H70;
		32'H00380001: READ <= 8'H70;
		32'H00380002: READ <= 8'H70;
		32'H00380003: READ <= 8'H6f;
		32'H00380004: READ <= 8'H6f;
		32'H00380005: READ <= 8'H6e;
		32'H00380006: READ <= 8'H6e;
		32'H00380007: READ <= 8'H6d;
		32'H00380008: READ <= 8'H6d;
		32'H00380009: READ <= 8'H6d;
		32'H0038000a: READ <= 8'H6d;
		32'H0038000b: READ <= 8'H6c;
		32'H0038000c: READ <= 8'H6c;
		32'H0038000d: READ <= 8'H6c;
		32'H0038000e: READ <= 8'H6c;
		32'H0038000f: READ <= 8'H6c;
		32'H00380010: READ <= 8'H6c;
		32'H00380011: READ <= 8'H6d;
		32'H00380012: READ <= 8'H6e;
		32'H00380013: READ <= 8'H6f;
		32'H00380014: READ <= 8'H72;
		32'H00380015: READ <= 8'H73;
		32'H00380016: READ <= 8'H74;
		32'H00380017: READ <= 8'H76;
		32'H00380018: READ <= 8'H78;
		32'H00380019: READ <= 8'H79;
		32'H0038001a: READ <= 8'H7c;
		32'H0038001b: READ <= 8'H7f;
		32'H0038001c: READ <= 8'H86;
		32'H0038001d: READ <= 8'H5b;
		32'H0038001e: READ <= 8'H64;
		32'H0038001f: READ <= 8'H79;
		32'H00380020: READ <= 8'H96;
		32'H00380021: READ <= 8'H8e;
		32'H00380022: READ <= 8'H8f;
		32'H00380023: READ <= 8'H74;
		32'H00380024: READ <= 8'H84;
		32'H00380025: READ <= 8'H46;
		32'H00380026: READ <= 8'H52;
		32'H00380027: READ <= 8'H52;
		32'H00380028: READ <= 8'H83;
		32'H00380029: READ <= 8'Hb7;
		32'H0038002a: READ <= 8'Hca;
		32'H0038002b: READ <= 8'Hd5;
		32'H0038002c: READ <= 8'Hdc;
		32'H0038002d: READ <= 8'Hdd;
		32'H0038002e: READ <= 8'Hde;
		32'H0038002f: READ <= 8'Hdf;
		32'H00380030: READ <= 8'He2;
		32'H00380031: READ <= 8'He2;
		32'H00380032: READ <= 8'He0;
		32'H00380033: READ <= 8'Hdd;
		32'H00380034: READ <= 8'Hda;
		32'H00380035: READ <= 8'Hd9;
		32'H00380036: READ <= 8'Hdc;
		32'H00380037: READ <= 8'Hde;
		32'H00380038: READ <= 8'He3;
		32'H00380039: READ <= 8'He3;
		32'H0038003a: READ <= 8'Hc1;
		32'H0038003b: READ <= 8'H6e;
		32'H0038003c: READ <= 8'H18;
		32'H0038003d: READ <= 8'H79;
		32'H0038003e: READ <= 8'H85;
		32'H0038003f: READ <= 8'H6f;
		32'H00380040: READ <= 8'H63;
		32'H00380041: READ <= 8'H77;
		32'H00380042: READ <= 8'H71;
		32'H00380043: READ <= 8'H75;
		32'H00380044: READ <= 8'H80;
		32'H00380045: READ <= 8'H91;
		32'H00380046: READ <= 8'H9b;
		32'H00380047: READ <= 8'Ha7;
		32'H00380048: READ <= 8'Haf;
		32'H00380049: READ <= 8'Ha3;
		32'H0038004a: READ <= 8'H8a;
		32'H0038004b: READ <= 8'H76;
		32'H0038004c: READ <= 8'H78;
		32'H0038004d: READ <= 8'H79;
		32'H0038004e: READ <= 8'H79;
		32'H0038004f: READ <= 8'H7a;
		32'H00380050: READ <= 8'H7a;
		32'H00380051: READ <= 8'H7b;
		32'H00380052: READ <= 8'H7c;
		32'H00380053: READ <= 8'H7d;
		32'H00380054: READ <= 8'H7e;
		32'H00380055: READ <= 8'H7e;
		32'H00380056: READ <= 8'H80;
		32'H00380057: READ <= 8'H80;
		32'H00380058: READ <= 8'H81;
		32'H00380059: READ <= 8'H82;
		32'H0038005a: READ <= 8'H83;
		32'H0038005b: READ <= 8'H84;
		32'H0038005c: READ <= 8'H86;
		32'H0038005d: READ <= 8'H87;
		32'H0038005e: READ <= 8'H88;
		32'H0038005f: READ <= 8'H88;
		32'H00380060: READ <= 8'H88;
		32'H00380061: READ <= 8'H89;
		32'H00380062: READ <= 8'H89;
		32'H00380063: READ <= 8'H89;
		
		32'H00390000: READ <= 8'H70;
		32'H00390001: READ <= 8'H70;
		32'H00390002: READ <= 8'H70;
		32'H00390003: READ <= 8'H6f;
		32'H00390004: READ <= 8'H6f;
		32'H00390005: READ <= 8'H6e;
		32'H00390006: READ <= 8'H6e;
		32'H00390007: READ <= 8'H6d;
		32'H00390008: READ <= 8'H6d;
		32'H00390009: READ <= 8'H6d;
		32'H0039000a: READ <= 8'H6c;
		32'H0039000b: READ <= 8'H6c;
		32'H0039000c: READ <= 8'H6b;
		32'H0039000d: READ <= 8'H6b;
		32'H0039000e: READ <= 8'H6b;
		32'H0039000f: READ <= 8'H6b;
		32'H00390010: READ <= 8'H6b;
		32'H00390011: READ <= 8'H6c;
		32'H00390012: READ <= 8'H6d;
		32'H00390013: READ <= 8'H6d;
		32'H00390014: READ <= 8'H6f;
		32'H00390015: READ <= 8'H71;
		32'H00390016: READ <= 8'H72;
		32'H00390017: READ <= 8'H73;
		32'H00390018: READ <= 8'H76;
		32'H00390019: READ <= 8'H77;
		32'H0039001a: READ <= 8'H7a;
		32'H0039001b: READ <= 8'H7e;
		32'H0039001c: READ <= 8'H80;
		32'H0039001d: READ <= 8'H87;
		32'H0039001e: READ <= 8'H8a;
		32'H0039001f: READ <= 8'H89;
		32'H00390020: READ <= 8'H87;
		32'H00390021: READ <= 8'H88;
		32'H00390022: READ <= 8'H8c;
		32'H00390023: READ <= 8'H96;
		32'H00390024: READ <= 8'H75;
		32'H00390025: READ <= 8'H5b;
		32'H00390026: READ <= 8'H6e;
		32'H00390027: READ <= 8'H65;
		32'H00390028: READ <= 8'H8f;
		32'H00390029: READ <= 8'Hbe;
		32'H0039002a: READ <= 8'Hcb;
		32'H0039002b: READ <= 8'Hd3;
		32'H0039002c: READ <= 8'Hd8;
		32'H0039002d: READ <= 8'Hd9;
		32'H0039002e: READ <= 8'Hd9;
		32'H0039002f: READ <= 8'Hda;
		32'H00390030: READ <= 8'Hdd;
		32'H00390031: READ <= 8'Hdd;
		32'H00390032: READ <= 8'Hdc;
		32'H00390033: READ <= 8'Hdc;
		32'H00390034: READ <= 8'Hdd;
		32'H00390035: READ <= 8'Hdf;
		32'H00390036: READ <= 8'He4;
		32'H00390037: READ <= 8'He5;
		32'H00390038: READ <= 8'He4;
		32'H00390039: READ <= 8'Hea;
		32'H0039003a: READ <= 8'He9;
		32'H0039003b: READ <= 8'H73;
		32'H0039003c: READ <= 8'H1b;
		32'H0039003d: READ <= 8'H73;
		32'H0039003e: READ <= 8'H8c;
		32'H0039003f: READ <= 8'H5f;
		32'H00390040: READ <= 8'H58;
		32'H00390041: READ <= 8'H74;
		32'H00390042: READ <= 8'H6e;
		32'H00390043: READ <= 8'H7f;
		32'H00390044: READ <= 8'H8d;
		32'H00390045: READ <= 8'H90;
		32'H00390046: READ <= 8'Ha5;
		32'H00390047: READ <= 8'Haf;
		32'H00390048: READ <= 8'Ha3;
		32'H00390049: READ <= 8'H96;
		32'H0039004a: READ <= 8'H79;
		32'H0039004b: READ <= 8'H77;
		32'H0039004c: READ <= 8'H78;
		32'H0039004d: READ <= 8'H78;
		32'H0039004e: READ <= 8'H79;
		32'H0039004f: READ <= 8'H7a;
		32'H00390050: READ <= 8'H7a;
		32'H00390051: READ <= 8'H7b;
		32'H00390052: READ <= 8'H7c;
		32'H00390053: READ <= 8'H7d;
		32'H00390054: READ <= 8'H7d;
		32'H00390055: READ <= 8'H7e;
		32'H00390056: READ <= 8'H7f;
		32'H00390057: READ <= 8'H80;
		32'H00390058: READ <= 8'H80;
		32'H00390059: READ <= 8'H82;
		32'H0039005a: READ <= 8'H83;
		32'H0039005b: READ <= 8'H85;
		32'H0039005c: READ <= 8'H86;
		32'H0039005d: READ <= 8'H86;
		32'H0039005e: READ <= 8'H87;
		32'H0039005f: READ <= 8'H88;
		32'H00390060: READ <= 8'H88;
		32'H00390061: READ <= 8'H88;
		32'H00390062: READ <= 8'H89;
		32'H00390063: READ <= 8'H8a;
		
		32'H003a0000: READ <= 8'H71;
		32'H003a0001: READ <= 8'H71;
		32'H003a0002: READ <= 8'H70;
		32'H003a0003: READ <= 8'H70;
		32'H003a0004: READ <= 8'H6f;
		32'H003a0005: READ <= 8'H6f;
		32'H003a0006: READ <= 8'H6e;
		32'H003a0007: READ <= 8'H6e;
		32'H003a0008: READ <= 8'H6d;
		32'H003a0009: READ <= 8'H6d;
		32'H003a000a: READ <= 8'H6c;
		32'H003a000b: READ <= 8'H6b;
		32'H003a000c: READ <= 8'H6b;
		32'H003a000d: READ <= 8'H6a;
		32'H003a000e: READ <= 8'H6b;
		32'H003a000f: READ <= 8'H6a;
		32'H003a0010: READ <= 8'H6a;
		32'H003a0011: READ <= 8'H6b;
		32'H003a0012: READ <= 8'H6b;
		32'H003a0013: READ <= 8'H6c;
		32'H003a0014: READ <= 8'H6d;
		32'H003a0015: READ <= 8'H6f;
		32'H003a0016: READ <= 8'H71;
		32'H003a0017: READ <= 8'H72;
		32'H003a0018: READ <= 8'H73;
		32'H003a0019: READ <= 8'H75;
		32'H003a001a: READ <= 8'H78;
		32'H003a001b: READ <= 8'H7c;
		32'H003a001c: READ <= 8'H7e;
		32'H003a001d: READ <= 8'H80;
		32'H003a001e: READ <= 8'H83;
		32'H003a001f: READ <= 8'H85;
		32'H003a0020: READ <= 8'H87;
		32'H003a0021: READ <= 8'H88;
		32'H003a0022: READ <= 8'H94;
		32'H003a0023: READ <= 8'H94;
		32'H003a0024: READ <= 8'H55;
		32'H003a0025: READ <= 8'H84;
		32'H003a0026: READ <= 8'H85;
		32'H003a0027: READ <= 8'H70;
		32'H003a0028: READ <= 8'H9c;
		32'H003a0029: READ <= 8'Hc9;
		32'H003a002a: READ <= 8'Hce;
		32'H003a002b: READ <= 8'Hd2;
		32'H003a002c: READ <= 8'Hd4;
		32'H003a002d: READ <= 8'Hd4;
		32'H003a002e: READ <= 8'Hd3;
		32'H003a002f: READ <= 8'Hd4;
		32'H003a0030: READ <= 8'Hd6;
		32'H003a0031: READ <= 8'Hd7;
		32'H003a0032: READ <= 8'Hd8;
		32'H003a0033: READ <= 8'Hdb;
		32'H003a0034: READ <= 8'Hdf;
		32'H003a0035: READ <= 8'He3;
		32'H003a0036: READ <= 8'He8;
		32'H003a0037: READ <= 8'He8;
		32'H003a0038: READ <= 8'He2;
		32'H003a0039: READ <= 8'He1;
		32'H003a003a: READ <= 8'He7;
		32'H003a003b: READ <= 8'H79;
		32'H003a003c: READ <= 8'H24;
		32'H003a003d: READ <= 8'H7f;
		32'H003a003e: READ <= 8'H8e;
		32'H003a003f: READ <= 8'H59;
		32'H003a0040: READ <= 8'H50;
		32'H003a0041: READ <= 8'H7f;
		32'H003a0042: READ <= 8'H7a;
		32'H003a0043: READ <= 8'H7e;
		32'H003a0044: READ <= 8'H8f;
		32'H003a0045: READ <= 8'H9a;
		32'H003a0046: READ <= 8'Ha8;
		32'H003a0047: READ <= 8'Ha6;
		32'H003a0048: READ <= 8'H98;
		32'H003a0049: READ <= 8'H7a;
		32'H003a004a: READ <= 8'H76;
		32'H003a004b: READ <= 8'H77;
		32'H003a004c: READ <= 8'H78;
		32'H003a004d: READ <= 8'H78;
		32'H003a004e: READ <= 8'H79;
		32'H003a004f: READ <= 8'H7a;
		32'H003a0050: READ <= 8'H7b;
		32'H003a0051: READ <= 8'H7b;
		32'H003a0052: READ <= 8'H7c;
		32'H003a0053: READ <= 8'H7c;
		32'H003a0054: READ <= 8'H7d;
		32'H003a0055: READ <= 8'H7e;
		32'H003a0056: READ <= 8'H7f;
		32'H003a0057: READ <= 8'H80;
		32'H003a0058: READ <= 8'H81;
		32'H003a0059: READ <= 8'H83;
		32'H003a005a: READ <= 8'H83;
		32'H003a005b: READ <= 8'H84;
		32'H003a005c: READ <= 8'H86;
		32'H003a005d: READ <= 8'H86;
		32'H003a005e: READ <= 8'H87;
		32'H003a005f: READ <= 8'H88;
		32'H003a0060: READ <= 8'H88;
		32'H003a0061: READ <= 8'H88;
		32'H003a0062: READ <= 8'H89;
		32'H003a0063: READ <= 8'H89;
		
		32'H003b0000: READ <= 8'H72;
		32'H003b0001: READ <= 8'H71;
		32'H003b0002: READ <= 8'H71;
		32'H003b0003: READ <= 8'H71;
		32'H003b0004: READ <= 8'H70;
		32'H003b0005: READ <= 8'H6f;
		32'H003b0006: READ <= 8'H6e;
		32'H003b0007: READ <= 8'H6e;
		32'H003b0008: READ <= 8'H6e;
		32'H003b0009: READ <= 8'H6d;
		32'H003b000a: READ <= 8'H6d;
		32'H003b000b: READ <= 8'H6b;
		32'H003b000c: READ <= 8'H6b;
		32'H003b000d: READ <= 8'H6a;
		32'H003b000e: READ <= 8'H6a;
		32'H003b000f: READ <= 8'H69;
		32'H003b0010: READ <= 8'H69;
		32'H003b0011: READ <= 8'H69;
		32'H003b0012: READ <= 8'H6a;
		32'H003b0013: READ <= 8'H6b;
		32'H003b0014: READ <= 8'H6c;
		32'H003b0015: READ <= 8'H6c;
		32'H003b0016: READ <= 8'H6e;
		32'H003b0017: READ <= 8'H71;
		32'H003b0018: READ <= 8'H72;
		32'H003b0019: READ <= 8'H74;
		32'H003b001a: READ <= 8'H76;
		32'H003b001b: READ <= 8'H7a;
		32'H003b001c: READ <= 8'H7d;
		32'H003b001d: READ <= 8'H80;
		32'H003b001e: READ <= 8'H83;
		32'H003b001f: READ <= 8'H87;
		32'H003b0020: READ <= 8'H8a;
		32'H003b0021: READ <= 8'H8c;
		32'H003b0022: READ <= 8'H9c;
		32'H003b0023: READ <= 8'H7e;
		32'H003b0024: READ <= 8'H5d;
		32'H003b0025: READ <= 8'H84;
		32'H003b0026: READ <= 8'H85;
		32'H003b0027: READ <= 8'H7a;
		32'H003b0028: READ <= 8'Hb4;
		32'H003b0029: READ <= 8'Hd6;
		32'H003b002a: READ <= 8'Hd2;
		32'H003b002b: READ <= 8'Hd0;
		32'H003b002c: READ <= 8'Hd0;
		32'H003b002d: READ <= 8'Hd0;
		32'H003b002e: READ <= 8'Hd1;
		32'H003b002f: READ <= 8'Hd1;
		32'H003b0030: READ <= 8'Hd2;
		32'H003b0031: READ <= 8'Hd3;
		32'H003b0032: READ <= 8'Hd6;
		32'H003b0033: READ <= 8'Hdb;
		32'H003b0034: READ <= 8'He0;
		32'H003b0035: READ <= 8'He5;
		32'H003b0036: READ <= 8'Hea;
		32'H003b0037: READ <= 8'Heb;
		32'H003b0038: READ <= 8'He6;
		32'H003b0039: READ <= 8'He5;
		32'H003b003a: READ <= 8'He4;
		32'H003b003b: READ <= 8'H98;
		32'H003b003c: READ <= 8'H27;
		32'H003b003d: READ <= 8'H7c;
		32'H003b003e: READ <= 8'H7d;
		32'H003b003f: READ <= 8'H5a;
		32'H003b0040: READ <= 8'H4c;
		32'H003b0041: READ <= 8'H89;
		32'H003b0042: READ <= 8'H72;
		32'H003b0043: READ <= 8'H90;
		32'H003b0044: READ <= 8'H95;
		32'H003b0045: READ <= 8'Ha3;
		32'H003b0046: READ <= 8'Ha0;
		32'H003b0047: READ <= 8'H98;
		32'H003b0048: READ <= 8'H8f;
		32'H003b0049: READ <= 8'H71;
		32'H003b004a: READ <= 8'H75;
		32'H003b004b: READ <= 8'H76;
		32'H003b004c: READ <= 8'H78;
		32'H003b004d: READ <= 8'H78;
		32'H003b004e: READ <= 8'H79;
		32'H003b004f: READ <= 8'H7a;
		32'H003b0050: READ <= 8'H7a;
		32'H003b0051: READ <= 8'H7b;
		32'H003b0052: READ <= 8'H7c;
		32'H003b0053: READ <= 8'H7c;
		32'H003b0054: READ <= 8'H7d;
		32'H003b0055: READ <= 8'H7e;
		32'H003b0056: READ <= 8'H7f;
		32'H003b0057: READ <= 8'H80;
		32'H003b0058: READ <= 8'H81;
		32'H003b0059: READ <= 8'H82;
		32'H003b005a: READ <= 8'H83;
		32'H003b005b: READ <= 8'H84;
		32'H003b005c: READ <= 8'H85;
		32'H003b005d: READ <= 8'H86;
		32'H003b005e: READ <= 8'H87;
		32'H003b005f: READ <= 8'H87;
		32'H003b0060: READ <= 8'H88;
		32'H003b0061: READ <= 8'H88;
		32'H003b0062: READ <= 8'H89;
		32'H003b0063: READ <= 8'H8a;
		
		32'H003c0000: READ <= 8'H71;
		32'H003c0001: READ <= 8'H71;
		32'H003c0002: READ <= 8'H71;
		32'H003c0003: READ <= 8'H71;
		32'H003c0004: READ <= 8'H70;
		32'H003c0005: READ <= 8'H70;
		32'H003c0006: READ <= 8'H6f;
		32'H003c0007: READ <= 8'H6e;
		32'H003c0008: READ <= 8'H6e;
		32'H003c0009: READ <= 8'H6d;
		32'H003c000a: READ <= 8'H6d;
		32'H003c000b: READ <= 8'H6c;
		32'H003c000c: READ <= 8'H6c;
		32'H003c000d: READ <= 8'H6b;
		32'H003c000e: READ <= 8'H6a;
		32'H003c000f: READ <= 8'H6a;
		32'H003c0010: READ <= 8'H69;
		32'H003c0011: READ <= 8'H69;
		32'H003c0012: READ <= 8'H68;
		32'H003c0013: READ <= 8'H68;
		32'H003c0014: READ <= 8'H6a;
		32'H003c0015: READ <= 8'H6a;
		32'H003c0016: READ <= 8'H6c;
		32'H003c0017: READ <= 8'H6e;
		32'H003c0018: READ <= 8'H70;
		32'H003c0019: READ <= 8'H73;
		32'H003c001a: READ <= 8'H76;
		32'H003c001b: READ <= 8'H79;
		32'H003c001c: READ <= 8'H7c;
		32'H003c001d: READ <= 8'H81;
		32'H003c001e: READ <= 8'H86;
		32'H003c001f: READ <= 8'H8a;
		32'H003c0020: READ <= 8'H8d;
		32'H003c0021: READ <= 8'H91;
		32'H003c0022: READ <= 8'H99;
		32'H003c0023: READ <= 8'H5a;
		32'H003c0024: READ <= 8'Ha6;
		32'H003c0025: READ <= 8'H8e;
		32'H003c0026: READ <= 8'H90;
		32'H003c0027: READ <= 8'H73;
		32'H003c0028: READ <= 8'Hca;
		32'H003c0029: READ <= 8'Hd9;
		32'H003c002a: READ <= 8'Hd4;
		32'H003c002b: READ <= 8'Hd1;
		32'H003c002c: READ <= 8'Hce;
		32'H003c002d: READ <= 8'Hce;
		32'H003c002e: READ <= 8'Hd1;
		32'H003c002f: READ <= 8'Hd0;
		32'H003c0030: READ <= 8'Hd0;
		32'H003c0031: READ <= 8'Hd1;
		32'H003c0032: READ <= 8'Hd5;
		32'H003c0033: READ <= 8'Hda;
		32'H003c0034: READ <= 8'Hde;
		32'H003c0035: READ <= 8'He4;
		32'H003c0036: READ <= 8'He9;
		32'H003c0037: READ <= 8'Heb;
		32'H003c0038: READ <= 8'He6;
		32'H003c0039: READ <= 8'Heb;
		32'H003c003a: READ <= 8'He7;
		32'H003c003b: READ <= 8'Hac;
		32'H003c003c: READ <= 8'H1b;
		32'H003c003d: READ <= 8'H63;
		32'H003c003e: READ <= 8'H6e;
		32'H003c003f: READ <= 8'H5a;
		32'H003c0040: READ <= 8'H47;
		32'H003c0041: READ <= 8'H7a;
		32'H003c0042: READ <= 8'H78;
		32'H003c0043: READ <= 8'H97;
		32'H003c0044: READ <= 8'H9d;
		32'H003c0045: READ <= 8'Ha7;
		32'H003c0046: READ <= 8'H9d;
		32'H003c0047: READ <= 8'H89;
		32'H003c0048: READ <= 8'H77;
		32'H003c0049: READ <= 8'H73;
		32'H003c004a: READ <= 8'H75;
		32'H003c004b: READ <= 8'H76;
		32'H003c004c: READ <= 8'H77;
		32'H003c004d: READ <= 8'H78;
		32'H003c004e: READ <= 8'H79;
		32'H003c004f: READ <= 8'H7a;
		32'H003c0050: READ <= 8'H7b;
		32'H003c0051: READ <= 8'H7b;
		32'H003c0052: READ <= 8'H7c;
		32'H003c0053: READ <= 8'H7d;
		32'H003c0054: READ <= 8'H7d;
		32'H003c0055: READ <= 8'H7e;
		32'H003c0056: READ <= 8'H7f;
		32'H003c0057: READ <= 8'H80;
		32'H003c0058: READ <= 8'H81;
		32'H003c0059: READ <= 8'H82;
		32'H003c005a: READ <= 8'H83;
		32'H003c005b: READ <= 8'H84;
		32'H003c005c: READ <= 8'H85;
		32'H003c005d: READ <= 8'H86;
		32'H003c005e: READ <= 8'H87;
		32'H003c005f: READ <= 8'H87;
		32'H003c0060: READ <= 8'H87;
		32'H003c0061: READ <= 8'H88;
		32'H003c0062: READ <= 8'H89;
		32'H003c0063: READ <= 8'H8a;
		
		32'H003d0000: READ <= 8'H72;
		32'H003d0001: READ <= 8'H72;
		32'H003d0002: READ <= 8'H71;
		32'H003d0003: READ <= 8'H71;
		32'H003d0004: READ <= 8'H70;
		32'H003d0005: READ <= 8'H6f;
		32'H003d0006: READ <= 8'H6f;
		32'H003d0007: READ <= 8'H6e;
		32'H003d0008: READ <= 8'H6e;
		32'H003d0009: READ <= 8'H6e;
		32'H003d000a: READ <= 8'H6d;
		32'H003d000b: READ <= 8'H6c;
		32'H003d000c: READ <= 8'H6c;
		32'H003d000d: READ <= 8'H6b;
		32'H003d000e: READ <= 8'H6a;
		32'H003d000f: READ <= 8'H6a;
		32'H003d0010: READ <= 8'H6a;
		32'H003d0011: READ <= 8'H69;
		32'H003d0012: READ <= 8'H69;
		32'H003d0013: READ <= 8'H69;
		32'H003d0014: READ <= 8'H68;
		32'H003d0015: READ <= 8'H69;
		32'H003d0016: READ <= 8'H6a;
		32'H003d0017: READ <= 8'H6c;
		32'H003d0018: READ <= 8'H6e;
		32'H003d0019: READ <= 8'H70;
		32'H003d001a: READ <= 8'H74;
		32'H003d001b: READ <= 8'H79;
		32'H003d001c: READ <= 8'H7e;
		32'H003d001d: READ <= 8'H83;
		32'H003d001e: READ <= 8'H89;
		32'H003d001f: READ <= 8'H8d;
		32'H003d0020: READ <= 8'H90;
		32'H003d0021: READ <= 8'H96;
		32'H003d0022: READ <= 8'H88;
		32'H003d0023: READ <= 8'H77;
		32'H003d0024: READ <= 8'Hc3;
		32'H003d0025: READ <= 8'Hbd;
		32'H003d0026: READ <= 8'Ha1;
		32'H003d0027: READ <= 8'H81;
		32'H003d0028: READ <= 8'Hce;
		32'H003d0029: READ <= 8'Hd8;
		32'H003d002a: READ <= 8'Hd4;
		32'H003d002b: READ <= 8'Hd0;
		32'H003d002c: READ <= 8'Hce;
		32'H003d002d: READ <= 8'Hce;
		32'H003d002e: READ <= 8'Hcf;
		32'H003d002f: READ <= 8'Hcf;
		32'H003d0030: READ <= 8'Hcf;
		32'H003d0031: READ <= 8'Hd1;
		32'H003d0032: READ <= 8'Hd5;
		32'H003d0033: READ <= 8'Hd9;
		32'H003d0034: READ <= 8'Hdd;
		32'H003d0035: READ <= 8'He2;
		32'H003d0036: READ <= 8'He7;
		32'H003d0037: READ <= 8'He9;
		32'H003d0038: READ <= 8'He7;
		32'H003d0039: READ <= 8'Hec;
		32'H003d003a: READ <= 8'He0;
		32'H003d003b: READ <= 8'Hb2;
		32'H003d003c: READ <= 8'H23;
		32'H003d003d: READ <= 8'H66;
		32'H003d003e: READ <= 8'H4b;
		32'H003d003f: READ <= 8'H5c;
		32'H003d0040: READ <= 8'H54;
		32'H003d0041: READ <= 8'H83;
		32'H003d0042: READ <= 8'H8b;
		32'H003d0043: READ <= 8'H9d;
		32'H003d0044: READ <= 8'H95;
		32'H003d0045: READ <= 8'H90;
		32'H003d0046: READ <= 8'H90;
		32'H003d0047: READ <= 8'H76;
		32'H003d0048: READ <= 8'H72;
		32'H003d0049: READ <= 8'H74;
		32'H003d004a: READ <= 8'H75;
		32'H003d004b: READ <= 8'H76;
		32'H003d004c: READ <= 8'H76;
		32'H003d004d: READ <= 8'H78;
		32'H003d004e: READ <= 8'H79;
		32'H003d004f: READ <= 8'H7a;
		32'H003d0050: READ <= 8'H7a;
		32'H003d0051: READ <= 8'H7b;
		32'H003d0052: READ <= 8'H7b;
		32'H003d0053: READ <= 8'H7d;
		32'H003d0054: READ <= 8'H7d;
		32'H003d0055: READ <= 8'H7e;
		32'H003d0056: READ <= 8'H7f;
		32'H003d0057: READ <= 8'H80;
		32'H003d0058: READ <= 8'H80;
		32'H003d0059: READ <= 8'H81;
		32'H003d005a: READ <= 8'H83;
		32'H003d005b: READ <= 8'H84;
		32'H003d005c: READ <= 8'H85;
		32'H003d005d: READ <= 8'H86;
		32'H003d005e: READ <= 8'H87;
		32'H003d005f: READ <= 8'H88;
		32'H003d0060: READ <= 8'H87;
		32'H003d0061: READ <= 8'H88;
		32'H003d0062: READ <= 8'H88;
		32'H003d0063: READ <= 8'H89;
		
		32'H003e0000: READ <= 8'H72;
		32'H003e0001: READ <= 8'H71;
		32'H003e0002: READ <= 8'H72;
		32'H003e0003: READ <= 8'H71;
		32'H003e0004: READ <= 8'H70;
		32'H003e0005: READ <= 8'H70;
		32'H003e0006: READ <= 8'H6f;
		32'H003e0007: READ <= 8'H6f;
		32'H003e0008: READ <= 8'H6f;
		32'H003e0009: READ <= 8'H6e;
		32'H003e000a: READ <= 8'H6e;
		32'H003e000b: READ <= 8'H6d;
		32'H003e000c: READ <= 8'H6d;
		32'H003e000d: READ <= 8'H6c;
		32'H003e000e: READ <= 8'H6b;
		32'H003e000f: READ <= 8'H6a;
		32'H003e0010: READ <= 8'H6a;
		32'H003e0011: READ <= 8'H6a;
		32'H003e0012: READ <= 8'H6a;
		32'H003e0013: READ <= 8'H69;
		32'H003e0014: READ <= 8'H69;
		32'H003e0015: READ <= 8'H69;
		32'H003e0016: READ <= 8'H6a;
		32'H003e0017: READ <= 8'H6b;
		32'H003e0018: READ <= 8'H6b;
		32'H003e0019: READ <= 8'H6e;
		32'H003e001a: READ <= 8'H72;
		32'H003e001b: READ <= 8'H79;
		32'H003e001c: READ <= 8'H80;
		32'H003e001d: READ <= 8'H85;
		32'H003e001e: READ <= 8'H8b;
		32'H003e001f: READ <= 8'H8f;
		32'H003e0020: READ <= 8'H93;
		32'H003e0021: READ <= 8'H9c;
		32'H003e0022: READ <= 8'H74;
		32'H003e0023: READ <= 8'H94;
		32'H003e0024: READ <= 8'Hae;
		32'H003e0025: READ <= 8'Hb6;
		32'H003e0026: READ <= 8'Ha0;
		32'H003e0027: READ <= 8'H80;
		32'H003e0028: READ <= 8'Hc9;
		32'H003e0029: READ <= 8'Hd7;
		32'H003e002a: READ <= 8'Hd2;
		32'H003e002b: READ <= 8'Hd0;
		32'H003e002c: READ <= 8'Hce;
		32'H003e002d: READ <= 8'Hcf;
		32'H003e002e: READ <= 8'Hcf;
		32'H003e002f: READ <= 8'Hcf;
		32'H003e0030: READ <= 8'Hcf;
		32'H003e0031: READ <= 8'Hd1;
		32'H003e0032: READ <= 8'Hd4;
		32'H003e0033: READ <= 8'Hd8;
		32'H003e0034: READ <= 8'Hda;
		32'H003e0035: READ <= 8'Hde;
		32'H003e0036: READ <= 8'He2;
		32'H003e0037: READ <= 8'He5;
		32'H003e0038: READ <= 8'He5;
		32'H003e0039: READ <= 8'Hec;
		32'H003e003a: READ <= 8'Hd6;
		32'H003e003b: READ <= 8'H9b;
		32'H003e003c: READ <= 8'H62;
		32'H003e003d: READ <= 8'H7f;
		32'H003e003e: READ <= 8'H58;
		32'H003e003f: READ <= 8'H49;
		32'H003e0040: READ <= 8'H5a;
		32'H003e0041: READ <= 8'H91;
		32'H003e0042: READ <= 8'H8c;
		32'H003e0043: READ <= 8'H8f;
		32'H003e0044: READ <= 8'H9e;
		32'H003e0045: READ <= 8'H8f;
		32'H003e0046: READ <= 8'H76;
		32'H003e0047: READ <= 8'H71;
		32'H003e0048: READ <= 8'H71;
		32'H003e0049: READ <= 8'H73;
		32'H003e004a: READ <= 8'H74;
		32'H003e004b: READ <= 8'H76;
		32'H003e004c: READ <= 8'H77;
		32'H003e004d: READ <= 8'H78;
		32'H003e004e: READ <= 8'H79;
		32'H003e004f: READ <= 8'H7a;
		32'H003e0050: READ <= 8'H7a;
		32'H003e0051: READ <= 8'H7b;
		32'H003e0052: READ <= 8'H7c;
		32'H003e0053: READ <= 8'H7c;
		32'H003e0054: READ <= 8'H7d;
		32'H003e0055: READ <= 8'H7e;
		32'H003e0056: READ <= 8'H7f;
		32'H003e0057: READ <= 8'H80;
		32'H003e0058: READ <= 8'H80;
		32'H003e0059: READ <= 8'H82;
		32'H003e005a: READ <= 8'H83;
		32'H003e005b: READ <= 8'H84;
		32'H003e005c: READ <= 8'H85;
		32'H003e005d: READ <= 8'H86;
		32'H003e005e: READ <= 8'H87;
		32'H003e005f: READ <= 8'H87;
		32'H003e0060: READ <= 8'H87;
		32'H003e0061: READ <= 8'H88;
		32'H003e0062: READ <= 8'H88;
		32'H003e0063: READ <= 8'H89;
		
		32'H003f0000: READ <= 8'H72;
		32'H003f0001: READ <= 8'H72;
		32'H003f0002: READ <= 8'H71;
		32'H003f0003: READ <= 8'H70;
		32'H003f0004: READ <= 8'H70;
		32'H003f0005: READ <= 8'H70;
		32'H003f0006: READ <= 8'H70;
		32'H003f0007: READ <= 8'H6f;
		32'H003f0008: READ <= 8'H6f;
		32'H003f0009: READ <= 8'H6f;
		32'H003f000a: READ <= 8'H6e;
		32'H003f000b: READ <= 8'H6e;
		32'H003f000c: READ <= 8'H6d;
		32'H003f000d: READ <= 8'H6c;
		32'H003f000e: READ <= 8'H6c;
		32'H003f000f: READ <= 8'H6b;
		32'H003f0010: READ <= 8'H6a;
		32'H003f0011: READ <= 8'H6a;
		32'H003f0012: READ <= 8'H6a;
		32'H003f0013: READ <= 8'H6a;
		32'H003f0014: READ <= 8'H6a;
		32'H003f0015: READ <= 8'H6a;
		32'H003f0016: READ <= 8'H6a;
		32'H003f0017: READ <= 8'H6b;
		32'H003f0018: READ <= 8'H6b;
		32'H003f0019: READ <= 8'H6e;
		32'H003f001a: READ <= 8'H72;
		32'H003f001b: READ <= 8'H79;
		32'H003f001c: READ <= 8'H81;
		32'H003f001d: READ <= 8'H88;
		32'H003f001e: READ <= 8'H8e;
		32'H003f001f: READ <= 8'H92;
		32'H003f0020: READ <= 8'H96;
		32'H003f0021: READ <= 8'H9a;
		32'H003f0022: READ <= 8'H81;
		32'H003f0023: READ <= 8'H96;
		32'H003f0024: READ <= 8'Hc0;
		32'H003f0025: READ <= 8'Hcb;
		32'H003f0026: READ <= 8'Hae;
		32'H003f0027: READ <= 8'H8d;
		32'H003f0028: READ <= 8'Hc4;
		32'H003f0029: READ <= 8'Hd3;
		32'H003f002a: READ <= 8'Hd0;
		32'H003f002b: READ <= 8'Hcf;
		32'H003f002c: READ <= 8'Hcd;
		32'H003f002d: READ <= 8'Hcf;
		32'H003f002e: READ <= 8'Hcf;
		32'H003f002f: READ <= 8'Hce;
		32'H003f0030: READ <= 8'Hce;
		32'H003f0031: READ <= 8'Hd0;
		32'H003f0032: READ <= 8'Hd3;
		32'H003f0033: READ <= 8'Hd6;
		32'H003f0034: READ <= 8'Hd8;
		32'H003f0035: READ <= 8'Hda;
		32'H003f0036: READ <= 8'Hdb;
		32'H003f0037: READ <= 8'Hdb;
		32'H003f0038: READ <= 8'He3;
		32'H003f0039: READ <= 8'He8;
		32'H003f003a: READ <= 8'Hd3;
		32'H003f003b: READ <= 8'H61;
		32'H003f003c: READ <= 8'H77;
		32'H003f003d: READ <= 8'H93;
		32'H003f003e: READ <= 8'H57;
		32'H003f003f: READ <= 8'H53;
		32'H003f0040: READ <= 8'H80;
		32'H003f0041: READ <= 8'H94;
		32'H003f0042: READ <= 8'H98;
		32'H003f0043: READ <= 8'H8f;
		32'H003f0044: READ <= 8'H7d;
		32'H003f0045: READ <= 8'H73;
		32'H003f0046: READ <= 8'H70;
		32'H003f0047: READ <= 8'H71;
		32'H003f0048: READ <= 8'H71;
		32'H003f0049: READ <= 8'H72;
		32'H003f004a: READ <= 8'H74;
		32'H003f004b: READ <= 8'H75;
		32'H003f004c: READ <= 8'H76;
		32'H003f004d: READ <= 8'H78;
		32'H003f004e: READ <= 8'H78;
		32'H003f004f: READ <= 8'H7a;
		32'H003f0050: READ <= 8'H7a;
		32'H003f0051: READ <= 8'H7b;
		32'H003f0052: READ <= 8'H7c;
		32'H003f0053: READ <= 8'H7c;
		32'H003f0054: READ <= 8'H7d;
		32'H003f0055: READ <= 8'H7e;
		32'H003f0056: READ <= 8'H7e;
		32'H003f0057: READ <= 8'H80;
		32'H003f0058: READ <= 8'H80;
		32'H003f0059: READ <= 8'H82;
		32'H003f005a: READ <= 8'H83;
		32'H003f005b: READ <= 8'H84;
		32'H003f005c: READ <= 8'H84;
		32'H003f005d: READ <= 8'H85;
		32'H003f005e: READ <= 8'H86;
		32'H003f005f: READ <= 8'H87;
		32'H003f0060: READ <= 8'H87;
		32'H003f0061: READ <= 8'H88;
		32'H003f0062: READ <= 8'H88;
		32'H003f0063: READ <= 8'H88;
		
		32'H00400000: READ <= 8'H72;
		32'H00400001: READ <= 8'H71;
		32'H00400002: READ <= 8'H72;
		32'H00400003: READ <= 8'H71;
		32'H00400004: READ <= 8'H71;
		32'H00400005: READ <= 8'H70;
		32'H00400006: READ <= 8'H70;
		32'H00400007: READ <= 8'H70;
		32'H00400008: READ <= 8'H70;
		32'H00400009: READ <= 8'H6f;
		32'H0040000a: READ <= 8'H6e;
		32'H0040000b: READ <= 8'H6e;
		32'H0040000c: READ <= 8'H6d;
		32'H0040000d: READ <= 8'H6d;
		32'H0040000e: READ <= 8'H6c;
		32'H0040000f: READ <= 8'H6c;
		32'H00400010: READ <= 8'H6b;
		32'H00400011: READ <= 8'H6b;
		32'H00400012: READ <= 8'H6b;
		32'H00400013: READ <= 8'H6b;
		32'H00400014: READ <= 8'H6b;
		32'H00400015: READ <= 8'H6b;
		32'H00400016: READ <= 8'H6b;
		32'H00400017: READ <= 8'H6b;
		32'H00400018: READ <= 8'H6b;
		32'H00400019: READ <= 8'H6e;
		32'H0040001a: READ <= 8'H73;
		32'H0040001b: READ <= 8'H7a;
		32'H0040001c: READ <= 8'H82;
		32'H0040001d: READ <= 8'H8a;
		32'H0040001e: READ <= 8'H90;
		32'H0040001f: READ <= 8'H94;
		32'H00400020: READ <= 8'H99;
		32'H00400021: READ <= 8'H92;
		32'H00400022: READ <= 8'H85;
		32'H00400023: READ <= 8'Hab;
		32'H00400024: READ <= 8'Hca;
		32'H00400025: READ <= 8'Hdb;
		32'H00400026: READ <= 8'Hc3;
		32'H00400027: READ <= 8'Ha3;
		32'H00400028: READ <= 8'Hbc;
		32'H00400029: READ <= 8'Hcd;
		32'H0040002a: READ <= 8'Hce;
		32'H0040002b: READ <= 8'Hcf;
		32'H0040002c: READ <= 8'Hcd;
		32'H0040002d: READ <= 8'Hce;
		32'H0040002e: READ <= 8'Hcf;
		32'H0040002f: READ <= 8'Hcd;
		32'H00400030: READ <= 8'Hcd;
		32'H00400031: READ <= 8'Hce;
		32'H00400032: READ <= 8'Hd1;
		32'H00400033: READ <= 8'Hd3;
		32'H00400034: READ <= 8'Hd6;
		32'H00400035: READ <= 8'Hd8;
		32'H00400036: READ <= 8'Hd6;
		32'H00400037: READ <= 8'Hcc;
		32'H00400038: READ <= 8'Hde;
		32'H00400039: READ <= 8'Hd6;
		32'H0040003a: READ <= 8'Haa;
		32'H0040003b: READ <= 8'H5a;
		32'H0040003c: READ <= 8'Ha4;
		32'H0040003d: READ <= 8'H9f;
		32'H0040003e: READ <= 8'H8e;
		32'H0040003f: READ <= 8'H91;
		32'H00400040: READ <= 8'Had;
		32'H00400041: READ <= 8'H91;
		32'H00400042: READ <= 8'H94;
		32'H00400043: READ <= 8'H7a;
		32'H00400044: READ <= 8'H78;
		32'H00400045: READ <= 8'H73;
		32'H00400046: READ <= 8'H71;
		32'H00400047: READ <= 8'H71;
		32'H00400048: READ <= 8'H72;
		32'H00400049: READ <= 8'H73;
		32'H0040004a: READ <= 8'H74;
		32'H0040004b: READ <= 8'H75;
		32'H0040004c: READ <= 8'H76;
		32'H0040004d: READ <= 8'H77;
		32'H0040004e: READ <= 8'H78;
		32'H0040004f: READ <= 8'H79;
		32'H00400050: READ <= 8'H7b;
		32'H00400051: READ <= 8'H7b;
		32'H00400052: READ <= 8'H7c;
		32'H00400053: READ <= 8'H7c;
		32'H00400054: READ <= 8'H7d;
		32'H00400055: READ <= 8'H7d;
		32'H00400056: READ <= 8'H7e;
		32'H00400057: READ <= 8'H7f;
		32'H00400058: READ <= 8'H80;
		32'H00400059: READ <= 8'H81;
		32'H0040005a: READ <= 8'H83;
		32'H0040005b: READ <= 8'H84;
		32'H0040005c: READ <= 8'H84;
		32'H0040005d: READ <= 8'H85;
		32'H0040005e: READ <= 8'H86;
		32'H0040005f: READ <= 8'H86;
		32'H00400060: READ <= 8'H87;
		32'H00400061: READ <= 8'H88;
		32'H00400062: READ <= 8'H88;
		32'H00400063: READ <= 8'H88;
		
		32'H00410000: READ <= 8'H73;
		32'H00410001: READ <= 8'H72;
		32'H00410002: READ <= 8'H72;
		32'H00410003: READ <= 8'H71;
		32'H00410004: READ <= 8'H71;
		32'H00410005: READ <= 8'H70;
		32'H00410006: READ <= 8'H70;
		32'H00410007: READ <= 8'H70;
		32'H00410008: READ <= 8'H70;
		32'H00410009: READ <= 8'H6f;
		32'H0041000a: READ <= 8'H6f;
		32'H0041000b: READ <= 8'H6f;
		32'H0041000c: READ <= 8'H6e;
		32'H0041000d: READ <= 8'H6d;
		32'H0041000e: READ <= 8'H6d;
		32'H0041000f: READ <= 8'H6d;
		32'H00410010: READ <= 8'H6c;
		32'H00410011: READ <= 8'H6c;
		32'H00410012: READ <= 8'H6c;
		32'H00410013: READ <= 8'H6b;
		32'H00410014: READ <= 8'H6c;
		32'H00410015: READ <= 8'H6b;
		32'H00410016: READ <= 8'H6c;
		32'H00410017: READ <= 8'H6c;
		32'H00410018: READ <= 8'H6c;
		32'H00410019: READ <= 8'H70;
		32'H0041001a: READ <= 8'H75;
		32'H0041001b: READ <= 8'H7c;
		32'H0041001c: READ <= 8'H85;
		32'H0041001d: READ <= 8'H8c;
		32'H0041001e: READ <= 8'H92;
		32'H0041001f: READ <= 8'H97;
		32'H00410020: READ <= 8'H99;
		32'H00410021: READ <= 8'H7f;
		32'H00410022: READ <= 8'H9a;
		32'H00410023: READ <= 8'Hd1;
		32'H00410024: READ <= 8'Hd0;
		32'H00410025: READ <= 8'Hdb;
		32'H00410026: READ <= 8'Hcd;
		32'H00410027: READ <= 8'Hb9;
		32'H00410028: READ <= 8'Hbc;
		32'H00410029: READ <= 8'Hc8;
		32'H0041002a: READ <= 8'Hcd;
		32'H0041002b: READ <= 8'Hd0;
		32'H0041002c: READ <= 8'Hce;
		32'H0041002d: READ <= 8'Hce;
		32'H0041002e: READ <= 8'Hcf;
		32'H0041002f: READ <= 8'Hcd;
		32'H00410030: READ <= 8'Hcc;
		32'H00410031: READ <= 8'Hcc;
		32'H00410032: READ <= 8'Hce;
		32'H00410033: READ <= 8'Hd0;
		32'H00410034: READ <= 8'Hd2;
		32'H00410035: READ <= 8'Hd5;
		32'H00410036: READ <= 8'Hd8;
		32'H00410037: READ <= 8'Hcf;
		32'H00410038: READ <= 8'Hdd;
		32'H00410039: READ <= 8'Hb5;
		32'H0041003a: READ <= 8'H68;
		32'H0041003b: READ <= 8'Ha2;
		32'H0041003c: READ <= 8'Hb5;
		32'H0041003d: READ <= 8'Ha9;
		32'H0041003e: READ <= 8'H9b;
		32'H0041003f: READ <= 8'H98;
		32'H00410040: READ <= 8'H87;
		32'H00410041: READ <= 8'H82;
		32'H00410042: READ <= 8'H7f;
		32'H00410043: READ <= 8'H7d;
		32'H00410044: READ <= 8'H78;
		32'H00410045: READ <= 8'H75;
		32'H00410046: READ <= 8'H72;
		32'H00410047: READ <= 8'H71;
		32'H00410048: READ <= 8'H71;
		32'H00410049: READ <= 8'H72;
		32'H0041004a: READ <= 8'H74;
		32'H0041004b: READ <= 8'H75;
		32'H0041004c: READ <= 8'H76;
		32'H0041004d: READ <= 8'H78;
		32'H0041004e: READ <= 8'H79;
		32'H0041004f: READ <= 8'H7a;
		32'H00410050: READ <= 8'H7a;
		32'H00410051: READ <= 8'H7a;
		32'H00410052: READ <= 8'H7b;
		32'H00410053: READ <= 8'H7c;
		32'H00410054: READ <= 8'H7d;
		32'H00410055: READ <= 8'H7d;
		32'H00410056: READ <= 8'H7e;
		32'H00410057: READ <= 8'H80;
		32'H00410058: READ <= 8'H80;
		32'H00410059: READ <= 8'H82;
		32'H0041005a: READ <= 8'H82;
		32'H0041005b: READ <= 8'H83;
		32'H0041005c: READ <= 8'H85;
		32'H0041005d: READ <= 8'H85;
		32'H0041005e: READ <= 8'H86;
		32'H0041005f: READ <= 8'H86;
		32'H00410060: READ <= 8'H86;
		32'H00410061: READ <= 8'H88;
		32'H00410062: READ <= 8'H88;
		32'H00410063: READ <= 8'H88;
		
		32'H00420000: READ <= 8'H73;
		32'H00420001: READ <= 8'H73;
		32'H00420002: READ <= 8'H73;
		32'H00420003: READ <= 8'H72;
		32'H00420004: READ <= 8'H72;
		32'H00420005: READ <= 8'H71;
		32'H00420006: READ <= 8'H70;
		32'H00420007: READ <= 8'H70;
		32'H00420008: READ <= 8'H70;
		32'H00420009: READ <= 8'H70;
		32'H0042000a: READ <= 8'H70;
		32'H0042000b: READ <= 8'H6f;
		32'H0042000c: READ <= 8'H6f;
		32'H0042000d: READ <= 8'H6f;
		32'H0042000e: READ <= 8'H6e;
		32'H0042000f: READ <= 8'H6d;
		32'H00420010: READ <= 8'H6c;
		32'H00420011: READ <= 8'H6d;
		32'H00420012: READ <= 8'H6d;
		32'H00420013: READ <= 8'H6c;
		32'H00420014: READ <= 8'H6c;
		32'H00420015: READ <= 8'H6c;
		32'H00420016: READ <= 8'H6c;
		32'H00420017: READ <= 8'H6c;
		32'H00420018: READ <= 8'H6e;
		32'H00420019: READ <= 8'H71;
		32'H0042001a: READ <= 8'H77;
		32'H0042001b: READ <= 8'H7e;
		32'H0042001c: READ <= 8'H87;
		32'H0042001d: READ <= 8'H8e;
		32'H0042001e: READ <= 8'H95;
		32'H0042001f: READ <= 8'H98;
		32'H00420020: READ <= 8'H98;
		32'H00420021: READ <= 8'H80;
		32'H00420022: READ <= 8'Ha0;
		32'H00420023: READ <= 8'Hdf;
		32'H00420024: READ <= 8'Hd9;
		32'H00420025: READ <= 8'Hd9;
		32'H00420026: READ <= 8'Hd4;
		32'H00420027: READ <= 8'Hc9;
		32'H00420028: READ <= 8'Hc4;
		32'H00420029: READ <= 8'Hc7;
		32'H0042002a: READ <= 8'Hcf;
		32'H0042002b: READ <= 8'Hd2;
		32'H0042002c: READ <= 8'Hd0;
		32'H0042002d: READ <= 8'Hcf;
		32'H0042002e: READ <= 8'Hcf;
		32'H0042002f: READ <= 8'Hce;
		32'H00420030: READ <= 8'Hcd;
		32'H00420031: READ <= 8'Hcc;
		32'H00420032: READ <= 8'Hcc;
		32'H00420033: READ <= 8'Hcc;
		32'H00420034: READ <= 8'Hcd;
		32'H00420035: READ <= 8'Hd0;
		32'H00420036: READ <= 8'Hda;
		32'H00420037: READ <= 8'Hdc;
		32'H00420038: READ <= 8'Hcd;
		32'H00420039: READ <= 8'Ha1;
		32'H0042003a: READ <= 8'H91;
		32'H0042003b: READ <= 8'Hc0;
		32'H0042003c: READ <= 8'Hba;
		32'H0042003d: READ <= 8'Hb1;
		32'H0042003e: READ <= 8'Ha4;
		32'H0042003f: READ <= 8'H97;
		32'H00420040: READ <= 8'H8f;
		32'H00420041: READ <= 8'H89;
		32'H00420042: READ <= 8'H84;
		32'H00420043: READ <= 8'H7f;
		32'H00420044: READ <= 8'H7c;
		32'H00420045: READ <= 8'H78;
		32'H00420046: READ <= 8'H75;
		32'H00420047: READ <= 8'H72;
		32'H00420048: READ <= 8'H72;
		32'H00420049: READ <= 8'H72;
		32'H0042004a: READ <= 8'H73;
		32'H0042004b: READ <= 8'H75;
		32'H0042004c: READ <= 8'H76;
		32'H0042004d: READ <= 8'H77;
		32'H0042004e: READ <= 8'H78;
		32'H0042004f: READ <= 8'H79;
		32'H00420050: READ <= 8'H7a;
		32'H00420051: READ <= 8'H7a;
		32'H00420052: READ <= 8'H7c;
		32'H00420053: READ <= 8'H7c;
		32'H00420054: READ <= 8'H7d;
		32'H00420055: READ <= 8'H7e;
		32'H00420056: READ <= 8'H7f;
		32'H00420057: READ <= 8'H7f;
		32'H00420058: READ <= 8'H81;
		32'H00420059: READ <= 8'H81;
		32'H0042005a: READ <= 8'H82;
		32'H0042005b: READ <= 8'H83;
		32'H0042005c: READ <= 8'H84;
		32'H0042005d: READ <= 8'H85;
		32'H0042005e: READ <= 8'H86;
		32'H0042005f: READ <= 8'H86;
		32'H00420060: READ <= 8'H86;
		32'H00420061: READ <= 8'H87;
		32'H00420062: READ <= 8'H88;
		32'H00420063: READ <= 8'H88;
		
		32'H00430000: READ <= 8'H73;
		32'H00430001: READ <= 8'H73;
		32'H00430002: READ <= 8'H73;
		32'H00430003: READ <= 8'H73;
		32'H00430004: READ <= 8'H72;
		32'H00430005: READ <= 8'H71;
		32'H00430006: READ <= 8'H70;
		32'H00430007: READ <= 8'H70;
		32'H00430008: READ <= 8'H70;
		32'H00430009: READ <= 8'H70;
		32'H0043000a: READ <= 8'H70;
		32'H0043000b: READ <= 8'H70;
		32'H0043000c: READ <= 8'H6f;
		32'H0043000d: READ <= 8'H6f;
		32'H0043000e: READ <= 8'H6e;
		32'H0043000f: READ <= 8'H6d;
		32'H00430010: READ <= 8'H6d;
		32'H00430011: READ <= 8'H6e;
		32'H00430012: READ <= 8'H6d;
		32'H00430013: READ <= 8'H6d;
		32'H00430014: READ <= 8'H6e;
		32'H00430015: READ <= 8'H6d;
		32'H00430016: READ <= 8'H6d;
		32'H00430017: READ <= 8'H6d;
		32'H00430018: READ <= 8'H6e;
		32'H00430019: READ <= 8'H73;
		32'H0043001a: READ <= 8'H79;
		32'H0043001b: READ <= 8'H7f;
		32'H0043001c: READ <= 8'H89;
		32'H0043001d: READ <= 8'H90;
		32'H0043001e: READ <= 8'H96;
		32'H0043001f: READ <= 8'H98;
		32'H00430020: READ <= 8'H9c;
		32'H00430021: READ <= 8'H7f;
		32'H00430022: READ <= 8'Ha9;
		32'H00430023: READ <= 8'He1;
		32'H00430024: READ <= 8'He1;
		32'H00430025: READ <= 8'Hdd;
		32'H00430026: READ <= 8'Hd8;
		32'H00430027: READ <= 8'Hd4;
		32'H00430028: READ <= 8'Hce;
		32'H00430029: READ <= 8'Hcd;
		32'H0043002a: READ <= 8'Hd1;
		32'H0043002b: READ <= 8'Hd4;
		32'H0043002c: READ <= 8'Hd3;
		32'H0043002d: READ <= 8'Hd1;
		32'H0043002e: READ <= 8'Hd0;
		32'H0043002f: READ <= 8'Hd0;
		32'H00430030: READ <= 8'Hce;
		32'H00430031: READ <= 8'Hcd;
		32'H00430032: READ <= 8'Hcb;
		32'H00430033: READ <= 8'Hca;
		32'H00430034: READ <= 8'Hc8;
		32'H00430035: READ <= 8'Hca;
		32'H00430036: READ <= 8'Hd7;
		32'H00430037: READ <= 8'He2;
		32'H00430038: READ <= 8'Hc7;
		32'H00430039: READ <= 8'H91;
		32'H0043003a: READ <= 8'Haf;
		32'H0043003b: READ <= 8'Hc5;
		32'H0043003c: READ <= 8'Hbf;
		32'H0043003d: READ <= 8'Hb7;
		32'H0043003e: READ <= 8'Hab;
		32'H0043003f: READ <= 8'H9d;
		32'H00430040: READ <= 8'H94;
		32'H00430041: READ <= 8'H8c;
		32'H00430042: READ <= 8'H87;
		32'H00430043: READ <= 8'H82;
		32'H00430044: READ <= 8'H7f;
		32'H00430045: READ <= 8'H7a;
		32'H00430046: READ <= 8'H77;
		32'H00430047: READ <= 8'H74;
		32'H00430048: READ <= 8'H73;
		32'H00430049: READ <= 8'H73;
		32'H0043004a: READ <= 8'H73;
		32'H0043004b: READ <= 8'H74;
		32'H0043004c: READ <= 8'H76;
		32'H0043004d: READ <= 8'H76;
		32'H0043004e: READ <= 8'H78;
		32'H0043004f: READ <= 8'H78;
		32'H00430050: READ <= 8'H7a;
		32'H00430051: READ <= 8'H7a;
		32'H00430052: READ <= 8'H7b;
		32'H00430053: READ <= 8'H7c;
		32'H00430054: READ <= 8'H7d;
		32'H00430055: READ <= 8'H7e;
		32'H00430056: READ <= 8'H7f;
		32'H00430057: READ <= 8'H7f;
		32'H00430058: READ <= 8'H81;
		32'H00430059: READ <= 8'H81;
		32'H0043005a: READ <= 8'H82;
		32'H0043005b: READ <= 8'H83;
		32'H0043005c: READ <= 8'H84;
		32'H0043005d: READ <= 8'H84;
		32'H0043005e: READ <= 8'H85;
		32'H0043005f: READ <= 8'H85;
		32'H00430060: READ <= 8'H86;
		32'H00430061: READ <= 8'H87;
		32'H00430062: READ <= 8'H88;
		32'H00430063: READ <= 8'H88;
		
		32'H00440000: READ <= 8'H74;
		32'H00440001: READ <= 8'H74;
		32'H00440002: READ <= 8'H74;
		32'H00440003: READ <= 8'H73;
		32'H00440004: READ <= 8'H72;
		32'H00440005: READ <= 8'H72;
		32'H00440006: READ <= 8'H71;
		32'H00440007: READ <= 8'H71;
		32'H00440008: READ <= 8'H70;
		32'H00440009: READ <= 8'H70;
		32'H0044000a: READ <= 8'H70;
		32'H0044000b: READ <= 8'H70;
		32'H0044000c: READ <= 8'H70;
		32'H0044000d: READ <= 8'H70;
		32'H0044000e: READ <= 8'H6f;
		32'H0044000f: READ <= 8'H6e;
		32'H00440010: READ <= 8'H6e;
		32'H00440011: READ <= 8'H6e;
		32'H00440012: READ <= 8'H6e;
		32'H00440013: READ <= 8'H6e;
		32'H00440014: READ <= 8'H6d;
		32'H00440015: READ <= 8'H6d;
		32'H00440016: READ <= 8'H6d;
		32'H00440017: READ <= 8'H6d;
		32'H00440018: READ <= 8'H6e;
		32'H00440019: READ <= 8'H74;
		32'H0044001a: READ <= 8'H7a;
		32'H0044001b: READ <= 8'H80;
		32'H0044001c: READ <= 8'H89;
		32'H0044001d: READ <= 8'H91;
		32'H0044001e: READ <= 8'H97;
		32'H0044001f: READ <= 8'H98;
		32'H00440020: READ <= 8'Ha8;
		32'H00440021: READ <= 8'H8e;
		32'H00440022: READ <= 8'Hcf;
		32'H00440023: READ <= 8'He5;
		32'H00440024: READ <= 8'He6;
		32'H00440025: READ <= 8'He4;
		32'H00440026: READ <= 8'Hdd;
		32'H00440027: READ <= 8'Hda;
		32'H00440028: READ <= 8'Hd8;
		32'H00440029: READ <= 8'Hd6;
		32'H0044002a: READ <= 8'Hd6;
		32'H0044002b: READ <= 8'Hd5;
		32'H0044002c: READ <= 8'Hd5;
		32'H0044002d: READ <= 8'Hd4;
		32'H0044002e: READ <= 8'Hd3;
		32'H0044002f: READ <= 8'Hd3;
		32'H00440030: READ <= 8'Hd1;
		32'H00440031: READ <= 8'Hcf;
		32'H00440032: READ <= 8'Hcd;
		32'H00440033: READ <= 8'Hcb;
		32'H00440034: READ <= 8'Hc6;
		32'H00440035: READ <= 8'Hc4;
		32'H00440036: READ <= 8'Hce;
		32'H00440037: READ <= 8'Hdc;
		32'H00440038: READ <= 8'Hce;
		32'H00440039: READ <= 8'H8b;
		32'H0044003a: READ <= 8'Hc8;
		32'H0044003b: READ <= 8'Hc9;
		32'H0044003c: READ <= 8'Hc3;
		32'H0044003d: READ <= 8'Hbb;
		32'H0044003e: READ <= 8'Hb0;
		32'H0044003f: READ <= 8'Ha3;
		32'H00440040: READ <= 8'H98;
		32'H00440041: READ <= 8'H91;
		32'H00440042: READ <= 8'H8a;
		32'H00440043: READ <= 8'H85;
		32'H00440044: READ <= 8'H81;
		32'H00440045: READ <= 8'H7d;
		32'H00440046: READ <= 8'H79;
		32'H00440047: READ <= 8'H77;
		32'H00440048: READ <= 8'H74;
		32'H00440049: READ <= 8'H73;
		32'H0044004a: READ <= 8'H73;
		32'H0044004b: READ <= 8'H75;
		32'H0044004c: READ <= 8'H76;
		32'H0044004d: READ <= 8'H76;
		32'H0044004e: READ <= 8'H78;
		32'H0044004f: READ <= 8'H79;
		32'H00440050: READ <= 8'H79;
		32'H00440051: READ <= 8'H7a;
		32'H00440052: READ <= 8'H7b;
		32'H00440053: READ <= 8'H7c;
		32'H00440054: READ <= 8'H7d;
		32'H00440055: READ <= 8'H7d;
		32'H00440056: READ <= 8'H7f;
		32'H00440057: READ <= 8'H80;
		32'H00440058: READ <= 8'H81;
		32'H00440059: READ <= 8'H81;
		32'H0044005a: READ <= 8'H82;
		32'H0044005b: READ <= 8'H83;
		32'H0044005c: READ <= 8'H84;
		32'H0044005d: READ <= 8'H84;
		32'H0044005e: READ <= 8'H85;
		32'H0044005f: READ <= 8'H86;
		32'H00440060: READ <= 8'H86;
		32'H00440061: READ <= 8'H87;
		32'H00440062: READ <= 8'H88;
		32'H00440063: READ <= 8'H88;
		
		32'H00450000: READ <= 8'H74;
		32'H00450001: READ <= 8'H74;
		32'H00450002: READ <= 8'H74;
		32'H00450003: READ <= 8'H74;
		32'H00450004: READ <= 8'H74;
		32'H00450005: READ <= 8'H73;
		32'H00450006: READ <= 8'H72;
		32'H00450007: READ <= 8'H72;
		32'H00450008: READ <= 8'H72;
		32'H00450009: READ <= 8'H71;
		32'H0045000a: READ <= 8'H71;
		32'H0045000b: READ <= 8'H70;
		32'H0045000c: READ <= 8'H70;
		32'H0045000d: READ <= 8'H70;
		32'H0045000e: READ <= 8'H6f;
		32'H0045000f: READ <= 8'H6f;
		32'H00450010: READ <= 8'H6f;
		32'H00450011: READ <= 8'H6f;
		32'H00450012: READ <= 8'H6e;
		32'H00450013: READ <= 8'H6e;
		32'H00450014: READ <= 8'H6e;
		32'H00450015: READ <= 8'H6e;
		32'H00450016: READ <= 8'H6d;
		32'H00450017: READ <= 8'H6e;
		32'H00450018: READ <= 8'H6f;
		32'H00450019: READ <= 8'H74;
		32'H0045001a: READ <= 8'H7b;
		32'H0045001b: READ <= 8'H82;
		32'H0045001c: READ <= 8'H8a;
		32'H0045001d: READ <= 8'H92;
		32'H0045001e: READ <= 8'H98;
		32'H0045001f: READ <= 8'H9b;
		32'H00450020: READ <= 8'Ha3;
		32'H00450021: READ <= 8'Hae;
		32'H00450022: READ <= 8'Hc7;
		32'H00450023: READ <= 8'Hde;
		32'H00450024: READ <= 8'He4;
		32'H00450025: READ <= 8'He4;
		32'H00450026: READ <= 8'Hdf;
		32'H00450027: READ <= 8'Hdd;
		32'H00450028: READ <= 8'Hdb;
		32'H00450029: READ <= 8'Hda;
		32'H0045002a: READ <= 8'Hd8;
		32'H0045002b: READ <= 8'Hd5;
		32'H0045002c: READ <= 8'Hd4;
		32'H0045002d: READ <= 8'Hd4;
		32'H0045002e: READ <= 8'Hd4;
		32'H0045002f: READ <= 8'Hd4;
		32'H00450030: READ <= 8'Hd1;
		32'H00450031: READ <= 8'Hce;
		32'H00450032: READ <= 8'Hcc;
		32'H00450033: READ <= 8'Hca;
		32'H00450034: READ <= 8'Hc7;
		32'H00450035: READ <= 8'Hc5;
		32'H00450036: READ <= 8'Hcc;
		32'H00450037: READ <= 8'Hdc;
		32'H00450038: READ <= 8'Ha3;
		32'H00450039: READ <= 8'Ha8;
		32'H0045003a: READ <= 8'Hd3;
		32'H0045003b: READ <= 8'Hcd;
		32'H0045003c: READ <= 8'Hc6;
		32'H0045003d: READ <= 8'Hbf;
		32'H0045003e: READ <= 8'Hb5;
		32'H0045003f: READ <= 8'Ha9;
		32'H00450040: READ <= 8'H9c;
		32'H00450041: READ <= 8'H94;
		32'H00450042: READ <= 8'H8e;
		32'H00450043: READ <= 8'H88;
		32'H00450044: READ <= 8'H84;
		32'H00450045: READ <= 8'H80;
		32'H00450046: READ <= 8'H7b;
		32'H00450047: READ <= 8'H78;
		32'H00450048: READ <= 8'H76;
		32'H00450049: READ <= 8'H73;
		32'H0045004a: READ <= 8'H73;
		32'H0045004b: READ <= 8'H74;
		32'H0045004c: READ <= 8'H75;
		32'H0045004d: READ <= 8'H76;
		32'H0045004e: READ <= 8'H77;
		32'H0045004f: READ <= 8'H78;
		32'H00450050: READ <= 8'H79;
		32'H00450051: READ <= 8'H7a;
		32'H00450052: READ <= 8'H7b;
		32'H00450053: READ <= 8'H7c;
		32'H00450054: READ <= 8'H7d;
		32'H00450055: READ <= 8'H7d;
		32'H00450056: READ <= 8'H7f;
		32'H00450057: READ <= 8'H7f;
		32'H00450058: READ <= 8'H80;
		32'H00450059: READ <= 8'H81;
		32'H0045005a: READ <= 8'H82;
		32'H0045005b: READ <= 8'H82;
		32'H0045005c: READ <= 8'H83;
		32'H0045005d: READ <= 8'H84;
		32'H0045005e: READ <= 8'H85;
		32'H0045005f: READ <= 8'H86;
		32'H00450060: READ <= 8'H86;
		32'H00450061: READ <= 8'H87;
		32'H00450062: READ <= 8'H88;
		32'H00450063: READ <= 8'H88;
		
		32'H00460000: READ <= 8'H74;
		32'H00460001: READ <= 8'H74;
		32'H00460002: READ <= 8'H74;
		32'H00460003: READ <= 8'H74;
		32'H00460004: READ <= 8'H74;
		32'H00460005: READ <= 8'H74;
		32'H00460006: READ <= 8'H73;
		32'H00460007: READ <= 8'H73;
		32'H00460008: READ <= 8'H73;
		32'H00460009: READ <= 8'H71;
		32'H0046000a: READ <= 8'H72;
		32'H0046000b: READ <= 8'H71;
		32'H0046000c: READ <= 8'H71;
		32'H0046000d: READ <= 8'H71;
		32'H0046000e: READ <= 8'H70;
		32'H0046000f: READ <= 8'H6f;
		32'H00460010: READ <= 8'H6f;
		32'H00460011: READ <= 8'H6f;
		32'H00460012: READ <= 8'H6f;
		32'H00460013: READ <= 8'H6f;
		32'H00460014: READ <= 8'H6e;
		32'H00460015: READ <= 8'H6e;
		32'H00460016: READ <= 8'H6e;
		32'H00460017: READ <= 8'H6e;
		32'H00460018: READ <= 8'H70;
		32'H00460019: READ <= 8'H75;
		32'H0046001a: READ <= 8'H7b;
		32'H0046001b: READ <= 8'H84;
		32'H0046001c: READ <= 8'H8b;
		32'H0046001d: READ <= 8'H92;
		32'H0046001e: READ <= 8'H99;
		32'H0046001f: READ <= 8'H9f;
		32'H00460020: READ <= 8'H9f;
		32'H00460021: READ <= 8'Hb9;
		32'H00460022: READ <= 8'Hb8;
		32'H00460023: READ <= 8'Hcd;
		32'H00460024: READ <= 8'Hdb;
		32'H00460025: READ <= 8'Hdf;
		32'H00460026: READ <= 8'Hde;
		32'H00460027: READ <= 8'Hdc;
		32'H00460028: READ <= 8'Hdc;
		32'H00460029: READ <= 8'Hdc;
		32'H0046002a: READ <= 8'Hda;
		32'H0046002b: READ <= 8'Hd6;
		32'H0046002c: READ <= 8'Hd4;
		32'H0046002d: READ <= 8'Hd4;
		32'H0046002e: READ <= 8'Hd3;
		32'H0046002f: READ <= 8'Hd2;
		32'H00460030: READ <= 8'Hd0;
		32'H00460031: READ <= 8'Hce;
		32'H00460032: READ <= 8'Hcd;
		32'H00460033: READ <= 8'Hca;
		32'H00460034: READ <= 8'Hc7;
		32'H00460035: READ <= 8'Hc8;
		32'H00460036: READ <= 8'Hce;
		32'H00460037: READ <= 8'Hbf;
		32'H00460038: READ <= 8'Haa;
		32'H00460039: READ <= 8'Hcd;
		32'H0046003a: READ <= 8'Hd5;
		32'H0046003b: READ <= 8'Hce;
		32'H0046003c: READ <= 8'Hca;
		32'H0046003d: READ <= 8'Hc3;
		32'H0046003e: READ <= 8'Hb9;
		32'H0046003f: READ <= 8'Had;
		32'H00460040: READ <= 8'Ha0;
		32'H00460041: READ <= 8'H97;
		32'H00460042: READ <= 8'H91;
		32'H00460043: READ <= 8'H8b;
		32'H00460044: READ <= 8'H86;
		32'H00460045: READ <= 8'H82;
		32'H00460046: READ <= 8'H7e;
		32'H00460047: READ <= 8'H7a;
		32'H00460048: READ <= 8'H78;
		32'H00460049: READ <= 8'H75;
		32'H0046004a: READ <= 8'H74;
		32'H0046004b: READ <= 8'H74;
		32'H0046004c: READ <= 8'H75;
		32'H0046004d: READ <= 8'H76;
		32'H0046004e: READ <= 8'H77;
		32'H0046004f: READ <= 8'H78;
		32'H00460050: READ <= 8'H79;
		32'H00460051: READ <= 8'H7a;
		32'H00460052: READ <= 8'H7b;
		32'H00460053: READ <= 8'H7c;
		32'H00460054: READ <= 8'H7d;
		32'H00460055: READ <= 8'H7d;
		32'H00460056: READ <= 8'H7e;
		32'H00460057: READ <= 8'H7f;
		32'H00460058: READ <= 8'H7f;
		32'H00460059: READ <= 8'H81;
		32'H0046005a: READ <= 8'H81;
		32'H0046005b: READ <= 8'H82;
		32'H0046005c: READ <= 8'H84;
		32'H0046005d: READ <= 8'H84;
		32'H0046005e: READ <= 8'H85;
		32'H0046005f: READ <= 8'H86;
		32'H00460060: READ <= 8'H86;
		32'H00460061: READ <= 8'H87;
		32'H00460062: READ <= 8'H87;
		32'H00460063: READ <= 8'H87;
		
		32'H00470000: READ <= 8'H75;
		32'H00470001: READ <= 8'H75;
		32'H00470002: READ <= 8'H75;
		32'H00470003: READ <= 8'H75;
		32'H00470004: READ <= 8'H75;
		32'H00470005: READ <= 8'H75;
		32'H00470006: READ <= 8'H74;
		32'H00470007: READ <= 8'H74;
		32'H00470008: READ <= 8'H73;
		32'H00470009: READ <= 8'H73;
		32'H0047000a: READ <= 8'H73;
		32'H0047000b: READ <= 8'H71;
		32'H0047000c: READ <= 8'H71;
		32'H0047000d: READ <= 8'H71;
		32'H0047000e: READ <= 8'H70;
		32'H0047000f: READ <= 8'H70;
		32'H00470010: READ <= 8'H70;
		32'H00470011: READ <= 8'H6f;
		32'H00470012: READ <= 8'H6f;
		32'H00470013: READ <= 8'H6f;
		32'H00470014: READ <= 8'H6f;
		32'H00470015: READ <= 8'H6e;
		32'H00470016: READ <= 8'H6f;
		32'H00470017: READ <= 8'H6f;
		32'H00470018: READ <= 8'H71;
		32'H00470019: READ <= 8'H76;
		32'H0047001a: READ <= 8'H7c;
		32'H0047001b: READ <= 8'H85;
		32'H0047001c: READ <= 8'H8e;
		32'H0047001d: READ <= 8'H94;
		32'H0047001e: READ <= 8'H9d;
		32'H0047001f: READ <= 8'Ha3;
		32'H00470020: READ <= 8'Hb5;
		32'H00470021: READ <= 8'Hba;
		32'H00470022: READ <= 8'Hb7;
		32'H00470023: READ <= 8'Hc1;
		32'H00470024: READ <= 8'Hd0;
		32'H00470025: READ <= 8'Hd9;
		32'H00470026: READ <= 8'Hda;
		32'H00470027: READ <= 8'Hdb;
		32'H00470028: READ <= 8'Hdc;
		32'H00470029: READ <= 8'Hdc;
		32'H0047002a: READ <= 8'Hdd;
		32'H0047002b: READ <= 8'Hd8;
		32'H0047002c: READ <= 8'Hd6;
		32'H0047002d: READ <= 8'Hd6;
		32'H0047002e: READ <= 8'Hd7;
		32'H0047002f: READ <= 8'Hd7;
		32'H00470030: READ <= 8'Hd6;
		32'H00470031: READ <= 8'Hd5;
		32'H00470032: READ <= 8'Hd2;
		32'H00470033: READ <= 8'Hd1;
		32'H00470034: READ <= 8'Hcf;
		32'H00470035: READ <= 8'Hd1;
		32'H00470036: READ <= 8'Hd6;
		32'H00470037: READ <= 8'Hd8;
		32'H00470038: READ <= 8'Hd7;
		32'H00470039: READ <= 8'Hd9;
		32'H0047003a: READ <= 8'Hd6;
		32'H0047003b: READ <= 8'Hd1;
		32'H0047003c: READ <= 8'Hcd;
		32'H0047003d: READ <= 8'Hc6;
		32'H0047003e: READ <= 8'Hbe;
		32'H0047003f: READ <= 8'Hb1;
		32'H00470040: READ <= 8'Ha4;
		32'H00470041: READ <= 8'H9b;
		32'H00470042: READ <= 8'H93;
		32'H00470043: READ <= 8'H8c;
		32'H00470044: READ <= 8'H88;
		32'H00470045: READ <= 8'H85;
		32'H00470046: READ <= 8'H80;
		32'H00470047: READ <= 8'H7b;
		32'H00470048: READ <= 8'H7a;
		32'H00470049: READ <= 8'H77;
		32'H0047004a: READ <= 8'H75;
		32'H0047004b: READ <= 8'H75;
		32'H0047004c: READ <= 8'H75;
		32'H0047004d: READ <= 8'H76;
		32'H0047004e: READ <= 8'H77;
		32'H0047004f: READ <= 8'H78;
		32'H00470050: READ <= 8'H79;
		32'H00470051: READ <= 8'H7a;
		32'H00470052: READ <= 8'H7b;
		32'H00470053: READ <= 8'H7b;
		32'H00470054: READ <= 8'H7d;
		32'H00470055: READ <= 8'H7d;
		32'H00470056: READ <= 8'H7e;
		32'H00470057: READ <= 8'H80;
		32'H00470058: READ <= 8'H7f;
		32'H00470059: READ <= 8'H81;
		32'H0047005a: READ <= 8'H82;
		32'H0047005b: READ <= 8'H82;
		32'H0047005c: READ <= 8'H82;
		32'H0047005d: READ <= 8'H84;
		32'H0047005e: READ <= 8'H85;
		32'H0047005f: READ <= 8'H86;
		32'H00470060: READ <= 8'H86;
		32'H00470061: READ <= 8'H86;
		32'H00470062: READ <= 8'H87;
		32'H00470063: READ <= 8'H87;
		
		32'H00480000: READ <= 8'H75;
		32'H00480001: READ <= 8'H76;
		32'H00480002: READ <= 8'H76;
		32'H00480003: READ <= 8'H75;
		32'H00480004: READ <= 8'H75;
		32'H00480005: READ <= 8'H75;
		32'H00480006: READ <= 8'H74;
		32'H00480007: READ <= 8'H75;
		32'H00480008: READ <= 8'H75;
		32'H00480009: READ <= 8'H74;
		32'H0048000a: READ <= 8'H73;
		32'H0048000b: READ <= 8'H73;
		32'H0048000c: READ <= 8'H72;
		32'H0048000d: READ <= 8'H71;
		32'H0048000e: READ <= 8'H71;
		32'H0048000f: READ <= 8'H71;
		32'H00480010: READ <= 8'H70;
		32'H00480011: READ <= 8'H70;
		32'H00480012: READ <= 8'H6f;
		32'H00480013: READ <= 8'H70;
		32'H00480014: READ <= 8'H6f;
		32'H00480015: READ <= 8'H6f;
		32'H00480016: READ <= 8'H6f;
		32'H00480017: READ <= 8'H70;
		32'H00480018: READ <= 8'H71;
		32'H00480019: READ <= 8'H77;
		32'H0048001a: READ <= 8'H7e;
		32'H0048001b: READ <= 8'H86;
		32'H0048001c: READ <= 8'H8f;
		32'H0048001d: READ <= 8'H97;
		32'H0048001e: READ <= 8'H9f;
		32'H0048001f: READ <= 8'Ha5;
		32'H00480020: READ <= 8'Hca;
		32'H00480021: READ <= 8'Hbd;
		32'H00480022: READ <= 8'Hb2;
		32'H00480023: READ <= 8'Hb7;
		32'H00480024: READ <= 8'Hc3;
		32'H00480025: READ <= 8'Hd0;
		32'H00480026: READ <= 8'Hd7;
		32'H00480027: READ <= 8'Hda;
		32'H00480028: READ <= 8'Hdc;
		32'H00480029: READ <= 8'Hdd;
		32'H0048002a: READ <= 8'Hde;
		32'H0048002b: READ <= 8'Hdb;
		32'H0048002c: READ <= 8'Hd9;
		32'H0048002d: READ <= 8'Hd8;
		32'H0048002e: READ <= 8'Hd9;
		32'H0048002f: READ <= 8'Hd9;
		32'H00480030: READ <= 8'Hd9;
		32'H00480031: READ <= 8'Hd8;
		32'H00480032: READ <= 8'Hd7;
		32'H00480033: READ <= 8'Hd6;
		32'H00480034: READ <= 8'Hd6;
		32'H00480035: READ <= 8'Hda;
		32'H00480036: READ <= 8'Hdb;
		32'H00480037: READ <= 8'Hdd;
		32'H00480038: READ <= 8'Hde;
		32'H00480039: READ <= 8'Hdb;
		32'H0048003a: READ <= 8'Hd7;
		32'H0048003b: READ <= 8'Hd3;
		32'H0048003c: READ <= 8'Hcf;
		32'H0048003d: READ <= 8'Hc9;
		32'H0048003e: READ <= 8'Hc0;
		32'H0048003f: READ <= 8'Hb5;
		32'H00480040: READ <= 8'Ha9;
		32'H00480041: READ <= 8'H9d;
		32'H00480042: READ <= 8'H96;
		32'H00480043: READ <= 8'H90;
		32'H00480044: READ <= 8'H8b;
		32'H00480045: READ <= 8'H87;
		32'H00480046: READ <= 8'H83;
		32'H00480047: READ <= 8'H7e;
		32'H00480048: READ <= 8'H7b;
		32'H00480049: READ <= 8'H78;
		32'H0048004a: READ <= 8'H76;
		32'H0048004b: READ <= 8'H76;
		32'H0048004c: READ <= 8'H75;
		32'H0048004d: READ <= 8'H75;
		32'H0048004e: READ <= 8'H77;
		32'H0048004f: READ <= 8'H78;
		32'H00480050: READ <= 8'H78;
		32'H00480051: READ <= 8'H79;
		32'H00480052: READ <= 8'H7b;
		32'H00480053: READ <= 8'H7b;
		32'H00480054: READ <= 8'H7c;
		32'H00480055: READ <= 8'H7c;
		32'H00480056: READ <= 8'H7e;
		32'H00480057: READ <= 8'H7f;
		32'H00480058: READ <= 8'H80;
		32'H00480059: READ <= 8'H81;
		32'H0048005a: READ <= 8'H82;
		32'H0048005b: READ <= 8'H82;
		32'H0048005c: READ <= 8'H83;
		32'H0048005d: READ <= 8'H84;
		32'H0048005e: READ <= 8'H85;
		32'H0048005f: READ <= 8'H85;
		32'H00480060: READ <= 8'H85;
		32'H00480061: READ <= 8'H86;
		32'H00480062: READ <= 8'H87;
		32'H00480063: READ <= 8'H87;
		
		32'H00490000: READ <= 8'H76;
		32'H00490001: READ <= 8'H76;
		32'H00490002: READ <= 8'H76;
		32'H00490003: READ <= 8'H76;
		32'H00490004: READ <= 8'H76;
		32'H00490005: READ <= 8'H76;
		32'H00490006: READ <= 8'H75;
		32'H00490007: READ <= 8'H75;
		32'H00490008: READ <= 8'H75;
		32'H00490009: READ <= 8'H74;
		32'H0049000a: READ <= 8'H74;
		32'H0049000b: READ <= 8'H74;
		32'H0049000c: READ <= 8'H73;
		32'H0049000d: READ <= 8'H72;
		32'H0049000e: READ <= 8'H73;
		32'H0049000f: READ <= 8'H71;
		32'H00490010: READ <= 8'H71;
		32'H00490011: READ <= 8'H70;
		32'H00490012: READ <= 8'H70;
		32'H00490013: READ <= 8'H70;
		32'H00490014: READ <= 8'H70;
		32'H00490015: READ <= 8'H70;
		32'H00490016: READ <= 8'H70;
		32'H00490017: READ <= 8'H70;
		32'H00490018: READ <= 8'H72;
		32'H00490019: READ <= 8'H77;
		32'H0049001a: READ <= 8'H7f;
		32'H0049001b: READ <= 8'H88;
		32'H0049001c: READ <= 8'H90;
		32'H0049001d: READ <= 8'H99;
		32'H0049001e: READ <= 8'Ha1;
		32'H0049001f: READ <= 8'Had;
		32'H00490020: READ <= 8'Hd0;
		32'H00490021: READ <= 8'Hb5;
		32'H00490022: READ <= 8'Ha0;
		32'H00490023: READ <= 8'Hb4;
		32'H00490024: READ <= 8'Hb6;
		32'H00490025: READ <= 8'Hc8;
		32'H00490026: READ <= 8'Hd3;
		32'H00490027: READ <= 8'Hd9;
		32'H00490028: READ <= 8'Hdb;
		32'H00490029: READ <= 8'Hdc;
		32'H0049002a: READ <= 8'Hde;
		32'H0049002b: READ <= 8'Hdd;
		32'H0049002c: READ <= 8'Hdc;
		32'H0049002d: READ <= 8'Hdc;
		32'H0049002e: READ <= 8'Hdd;
		32'H0049002f: READ <= 8'Hdd;
		32'H00490030: READ <= 8'Hdb;
		32'H00490031: READ <= 8'Hdb;
		32'H00490032: READ <= 8'Hdb;
		32'H00490033: READ <= 8'Hdc;
		32'H00490034: READ <= 8'Hdc;
		32'H00490035: READ <= 8'Hde;
		32'H00490036: READ <= 8'Hde;
		32'H00490037: READ <= 8'Hdf;
		32'H00490038: READ <= 8'He0;
		32'H00490039: READ <= 8'Hdd;
		32'H0049003a: READ <= 8'Hd9;
		32'H0049003b: READ <= 8'Hd5;
		32'H0049003c: READ <= 8'Hd0;
		32'H0049003d: READ <= 8'Hcc;
		32'H0049003e: READ <= 8'Hc4;
		32'H0049003f: READ <= 8'Hb9;
		32'H00490040: READ <= 8'Hac;
		32'H00490041: READ <= 8'Ha1;
		32'H00490042: READ <= 8'H99;
		32'H00490043: READ <= 8'H92;
		32'H00490044: READ <= 8'H8e;
		32'H00490045: READ <= 8'H89;
		32'H00490046: READ <= 8'H85;
		32'H00490047: READ <= 8'H80;
		32'H00490048: READ <= 8'H7d;
		32'H00490049: READ <= 8'H7a;
		32'H0049004a: READ <= 8'H77;
		32'H0049004b: READ <= 8'H78;
		32'H0049004c: READ <= 8'H76;
		32'H0049004d: READ <= 8'H76;
		32'H0049004e: READ <= 8'H77;
		32'H0049004f: READ <= 8'H78;
		32'H00490050: READ <= 8'H79;
		32'H00490051: READ <= 8'H79;
		32'H00490052: READ <= 8'H7b;
		32'H00490053: READ <= 8'H7b;
		32'H00490054: READ <= 8'H7c;
		32'H00490055: READ <= 8'H7d;
		32'H00490056: READ <= 8'H7e;
		32'H00490057: READ <= 8'H7e;
		32'H00490058: READ <= 8'H80;
		32'H00490059: READ <= 8'H80;
		32'H0049005a: READ <= 8'H81;
		32'H0049005b: READ <= 8'H83;
		32'H0049005c: READ <= 8'H83;
		32'H0049005d: READ <= 8'H83;
		32'H0049005e: READ <= 8'H85;
		32'H0049005f: READ <= 8'H85;
		32'H00490060: READ <= 8'H86;
		32'H00490061: READ <= 8'H86;
		32'H00490062: READ <= 8'H87;
		32'H00490063: READ <= 8'H86;
		
		32'H004a0000: READ <= 8'H76;
		32'H004a0001: READ <= 8'H76;
		32'H004a0002: READ <= 8'H76;
		32'H004a0003: READ <= 8'H75;
		32'H004a0004: READ <= 8'H76;
		32'H004a0005: READ <= 8'H76;
		32'H004a0006: READ <= 8'H76;
		32'H004a0007: READ <= 8'H75;
		32'H004a0008: READ <= 8'H76;
		32'H004a0009: READ <= 8'H75;
		32'H004a000a: READ <= 8'H74;
		32'H004a000b: READ <= 8'H74;
		32'H004a000c: READ <= 8'H74;
		32'H004a000d: READ <= 8'H73;
		32'H004a000e: READ <= 8'H73;
		32'H004a000f: READ <= 8'H71;
		32'H004a0010: READ <= 8'H71;
		32'H004a0011: READ <= 8'H71;
		32'H004a0012: READ <= 8'H70;
		32'H004a0013: READ <= 8'H70;
		32'H004a0014: READ <= 8'H70;
		32'H004a0015: READ <= 8'H70;
		32'H004a0016: READ <= 8'H70;
		32'H004a0017: READ <= 8'H71;
		32'H004a0018: READ <= 8'H74;
		32'H004a0019: READ <= 8'H78;
		32'H004a001a: READ <= 8'H7f;
		32'H004a001b: READ <= 8'H88;
		32'H004a001c: READ <= 8'H91;
		32'H004a001d: READ <= 8'H9b;
		32'H004a001e: READ <= 8'Ha3;
		32'H004a001f: READ <= 8'Hb6;
		32'H004a0020: READ <= 8'Hcd;
		32'H004a0021: READ <= 8'Hb5;
		32'H004a0022: READ <= 8'H9c;
		32'H004a0023: READ <= 8'Hab;
		32'H004a0024: READ <= 8'Hb6;
		32'H004a0025: READ <= 8'Hc3;
		32'H004a0026: READ <= 8'Hce;
		32'H004a0027: READ <= 8'Hd7;
		32'H004a0028: READ <= 8'Hda;
		32'H004a0029: READ <= 8'Hdc;
		32'H004a002a: READ <= 8'Hde;
		32'H004a002b: READ <= 8'Hdd;
		32'H004a002c: READ <= 8'Hdc;
		32'H004a002d: READ <= 8'Hdd;
		32'H004a002e: READ <= 8'Hde;
		32'H004a002f: READ <= 8'Hdf;
		32'H004a0030: READ <= 8'Hde;
		32'H004a0031: READ <= 8'Hde;
		32'H004a0032: READ <= 8'Hde;
		32'H004a0033: READ <= 8'Hdf;
		32'H004a0034: READ <= 8'Hdf;
		32'H004a0035: READ <= 8'He0;
		32'H004a0036: READ <= 8'He1;
		32'H004a0037: READ <= 8'He2;
		32'H004a0038: READ <= 8'He1;
		32'H004a0039: READ <= 8'Hde;
		32'H004a003a: READ <= 8'Hdb;
		32'H004a003b: READ <= 8'Hd6;
		32'H004a003c: READ <= 8'Hd2;
		32'H004a003d: READ <= 8'Hcd;
		32'H004a003e: READ <= 8'Hc6;
		32'H004a003f: READ <= 8'Hbb;
		32'H004a0040: READ <= 8'Hb0;
		32'H004a0041: READ <= 8'Ha4;
		32'H004a0042: READ <= 8'H9b;
		32'H004a0043: READ <= 8'H93;
		32'H004a0044: READ <= 8'H8f;
		32'H004a0045: READ <= 8'H8b;
		32'H004a0046: READ <= 8'H87;
		32'H004a0047: READ <= 8'H82;
		32'H004a0048: READ <= 8'H7f;
		32'H004a0049: READ <= 8'H7d;
		32'H004a004a: READ <= 8'H7a;
		32'H004a004b: READ <= 8'H77;
		32'H004a004c: READ <= 8'H76;
		32'H004a004d: READ <= 8'H77;
		32'H004a004e: READ <= 8'H77;
		32'H004a004f: READ <= 8'H77;
		32'H004a0050: READ <= 8'H78;
		32'H004a0051: READ <= 8'H79;
		32'H004a0052: READ <= 8'H7b;
		32'H004a0053: READ <= 8'H7c;
		32'H004a0054: READ <= 8'H7c;
		32'H004a0055: READ <= 8'H7d;
		32'H004a0056: READ <= 8'H7e;
		32'H004a0057: READ <= 8'H7e;
		32'H004a0058: READ <= 8'H7f;
		32'H004a0059: READ <= 8'H81;
		32'H004a005a: READ <= 8'H81;
		32'H004a005b: READ <= 8'H82;
		32'H004a005c: READ <= 8'H83;
		32'H004a005d: READ <= 8'H83;
		32'H004a005e: READ <= 8'H85;
		32'H004a005f: READ <= 8'H85;
		32'H004a0060: READ <= 8'H85;
		32'H004a0061: READ <= 8'H86;
		32'H004a0062: READ <= 8'H86;
		32'H004a0063: READ <= 8'H86;
		default: READ <= 8'b0;
	endcase
	end

endmodule
