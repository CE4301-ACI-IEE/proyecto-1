`timescale 1ns / 1ps
module mem_pic #( parameter SIZE = 8 )
(
  input logic CLK,
  input logic [SIZE-1:0] ADDRESS,
  output logic [SIZE-1:0] READ
);
always_ff@( posedge CLK ) begin
  case( ADDRESS << 2 )
      32'H0: READ <= 8'Hb3;
      32'H1: READ <= 8'Hb6;
      32'H2: READ <= 8'Hb8;
      32'H3: READ <= 8'Hbb;
      32'H4: READ <= 8'Hbe;
      32'H5: READ <= 8'Hc1;
      32'H6: READ <= 8'Hc5;
      32'H7: READ <= 8'Hc8;
      32'H8: READ <= 8'Hcb;
      32'H9: READ <= 8'Hce;
      32'H10: READ <= 8'Hd2;
      32'H11: READ <= 8'Hd5;
      32'H12: READ <= 8'Hd6;
      32'H13: READ <= 8'Hda;
      32'H14: READ <= 8'Hdc;
      32'H15: READ <= 8'Hdf;
      32'H16: READ <= 8'He1;
      32'H17: READ <= 8'He4;
      32'H18: READ <= 8'He6;
      32'H19: READ <= 8'He8;
      32'H20: READ <= 8'He9;
      32'H21: READ <= 8'Hea;
      32'H22: READ <= 8'Heb;
      32'H23: READ <= 8'Hec;
      32'H24: READ <= 8'Hee;
      32'H25: READ <= 8'Hee;
      32'H26: READ <= 8'Hef;
      32'H27: READ <= 8'Hef;
      32'H28: READ <= 8'Hf0;
      32'H29: READ <= 8'Hf1;
      32'H30: READ <= 8'Hf2;
      32'H31: READ <= 8'Hf2;
      32'H32: READ <= 8'Hf2;
      32'H33: READ <= 8'Hf2;
      32'H34: READ <= 8'Hf1;
      32'H35: READ <= 8'Hf0;
      32'H36: READ <= 8'Hef;
      32'H37: READ <= 8'Hee;
      32'H38: READ <= 8'Hed;
      32'H39: READ <= 8'Hea;
      32'H40: READ <= 8'He9;
      32'H41: READ <= 8'He8;
      32'H42: READ <= 8'He6;
      32'H43: READ <= 8'He2;
      32'H44: READ <= 8'He0;
      32'H45: READ <= 8'Hdc;
      32'H46: READ <= 8'Hd7;
      32'H47: READ <= 8'Hd3;
      32'H48: READ <= 8'Hce;
      32'H49: READ <= 8'Hc9;
      32'H50: READ <= 8'Hc3;
      32'H51: READ <= 8'Hbc;
      32'H52: READ <= 8'Hb3;
      32'H53: READ <= 8'Hac;
      32'H54: READ <= 8'Ha6;
      32'H55: READ <= 8'Ha1;
      32'H56: READ <= 8'H9f;
      32'H57: READ <= 8'H9d;
      32'H58: READ <= 8'H9c;
      32'H59: READ <= 8'H9b;
      32'H60: READ <= 8'H9b;
      32'H61: READ <= 8'H9b;
      32'H62: READ <= 8'H9a;
      32'H63: READ <= 8'H9b;
      32'H64: READ <= 8'H9b;
      32'H65: READ <= 8'H9b;
      32'H66: READ <= 8'H9c;
      32'H67: READ <= 8'H9d;
      32'H68: READ <= 8'H9d;
      32'H69: READ <= 8'H9d;
      32'H70: READ <= 8'H9d;
      32'H71: READ <= 8'H9d;
      32'H72: READ <= 8'H9e;
      32'H73: READ <= 8'H9d;
      32'H74: READ <= 8'H9e;
      32'H75: READ <= 8'H9f;
      32'H76: READ <= 8'H9f;
      32'H77: READ <= 8'H9f;
      32'H78: READ <= 8'Ha0;
      32'H79: READ <= 8'Ha1;
      32'H80: READ <= 8'Ha1;
      32'H81: READ <= 8'Ha2;
      32'H82: READ <= 8'Ha2;
      32'H83: READ <= 8'Ha3;
      32'H84: READ <= 8'Ha3;
      32'H85: READ <= 8'Ha3;
      32'H86: READ <= 8'Ha4;
      32'H87: READ <= 8'Ha4;
      32'H88: READ <= 8'Ha4;
      32'H89: READ <= 8'Ha4;
      32'H90: READ <= 8'Ha4;
      32'H91: READ <= 8'Ha3;
      32'H92: READ <= 8'Ha4;
      32'H93: READ <= 8'Ha4;
      32'H94: READ <= 8'Ha5;
      32'H95: READ <= 8'Ha5;
      32'H96: READ <= 8'Ha6;
      32'H97: READ <= 8'Ha7;
      32'H98: READ <= 8'Ha7;
      32'H99: READ <= 8'Ha8;
      32'H100: READ <= 8'Hb3;
      32'H101: READ <= 8'Hb5;
      32'H102: READ <= 8'Hb7;
      32'H103: READ <= 8'Hb9;
      32'H104: READ <= 8'Hbc;
      32'H105: READ <= 8'Hbf;
      32'H106: READ <= 8'Hc3;
      32'H107: READ <= 8'Hc6;
      32'H108: READ <= 8'Hc9;
      32'H109: READ <= 8'Hcd;
      32'H110: READ <= 8'Hd1;
      32'H111: READ <= 8'Hd3;
      32'H112: READ <= 8'Hd6;
      32'H113: READ <= 8'Hd9;
      32'H114: READ <= 8'Hdb;
      32'H115: READ <= 8'Hde;
      32'H116: READ <= 8'He0;
      32'H117: READ <= 8'He4;
      32'H118: READ <= 8'He6;
      32'H119: READ <= 8'He8;
      32'H120: READ <= 8'He9;
      32'H121: READ <= 8'Hea;
      32'H122: READ <= 8'Hec;
      32'H123: READ <= 8'Hec;
      32'H124: READ <= 8'Hee;
      32'H125: READ <= 8'Hee;
      32'H126: READ <= 8'Hef;
      32'H127: READ <= 8'Hf0;
      32'H128: READ <= 8'Hf0;
      32'H129: READ <= 8'Hf2;
      32'H130: READ <= 8'Hf2;
      32'H131: READ <= 8'Hf2;
      32'H132: READ <= 8'Hf2;
      32'H133: READ <= 8'Hf2;
      32'H134: READ <= 8'Hf2;
      32'H135: READ <= 8'Hf0;
      32'H136: READ <= 8'Hef;
      32'H137: READ <= 8'Hee;
      32'H138: READ <= 8'Hec;
      32'H139: READ <= 8'Heb;
      32'H140: READ <= 8'He9;
      32'H141: READ <= 8'He9;
      32'H142: READ <= 8'He7;
      32'H143: READ <= 8'He3;
      32'H144: READ <= 8'He0;
      32'H145: READ <= 8'Hdc;
      32'H146: READ <= 8'Hd8;
      32'H147: READ <= 8'Hd4;
      32'H148: READ <= 8'Hd0;
      32'H149: READ <= 8'Hcb;
      32'H150: READ <= 8'Hc5;
      32'H151: READ <= 8'Hbd;
      32'H152: READ <= 8'Hb4;
      32'H153: READ <= 8'Had;
      32'H154: READ <= 8'Ha6;
      32'H155: READ <= 8'Ha1;
      32'H156: READ <= 8'H9e;
      32'H157: READ <= 8'H9c;
      32'H158: READ <= 8'H9b;
      32'H159: READ <= 8'H9a;
      32'H160: READ <= 8'H9b;
      32'H161: READ <= 8'H9a;
      32'H162: READ <= 8'H99;
      32'H163: READ <= 8'H99;
      32'H164: READ <= 8'H9a;
      32'H165: READ <= 8'H9b;
      32'H166: READ <= 8'H9a;
      32'H167: READ <= 8'H9b;
      32'H168: READ <= 8'H9c;
      32'H169: READ <= 8'H9c;
      32'H170: READ <= 8'H9d;
      32'H171: READ <= 8'H9c;
      32'H172: READ <= 8'H9c;
      32'H173: READ <= 8'H9c;
      32'H174: READ <= 8'H9c;
      32'H175: READ <= 8'H9d;
      32'H176: READ <= 8'H9e;
      32'H177: READ <= 8'H9e;
      32'H178: READ <= 8'Ha0;
      32'H179: READ <= 8'Ha0;
      32'H180: READ <= 8'Ha0;
      32'H181: READ <= 8'Ha1;
      32'H182: READ <= 8'Ha1;
      32'H183: READ <= 8'Ha2;
      32'H184: READ <= 8'Ha3;
      32'H185: READ <= 8'Ha3;
      32'H186: READ <= 8'Ha2;
      32'H187: READ <= 8'Ha3;
      32'H188: READ <= 8'Ha3;
      32'H189: READ <= 8'Ha3;
      32'H190: READ <= 8'Ha3;
      32'H191: READ <= 8'Ha3;
      32'H192: READ <= 8'Ha3;
      32'H193: READ <= 8'Ha3;
      32'H194: READ <= 8'Ha4;
      32'H195: READ <= 8'Ha4;
      32'H196: READ <= 8'Ha6;
      32'H197: READ <= 8'Ha6;
      32'H198: READ <= 8'Ha6;
      32'H199: READ <= 8'Ha6;
      32'H200: READ <= 8'Hb1;
      32'H201: READ <= 8'Hb3;
      32'H202: READ <= 8'Hb6;
      32'H203: READ <= 8'Hb8;
      32'H204: READ <= 8'Hba;
      32'H205: READ <= 8'Hbd;
      32'H206: READ <= 8'Hc1;
      32'H207: READ <= 8'Hc5;
      32'H208: READ <= 8'Hc8;
      32'H209: READ <= 8'Hcc;
      32'H210: READ <= 8'Hcf;
      32'H211: READ <= 8'Hd2;
      32'H212: READ <= 8'Hd5;
      32'H213: READ <= 8'Hd8;
      32'H214: READ <= 8'Hda;
      32'H215: READ <= 8'Hdd;
      32'H216: READ <= 8'He0;
      32'H217: READ <= 8'He3;
      32'H218: READ <= 8'He5;
      32'H219: READ <= 8'He7;
      32'H220: READ <= 8'He9;
      32'H221: READ <= 8'Hea;
      32'H222: READ <= 8'Heb;
      32'H223: READ <= 8'Hec;
      32'H224: READ <= 8'Hee;
      32'H225: READ <= 8'Hee;
      32'H226: READ <= 8'Hef;
      32'H227: READ <= 8'Hef;
      32'H228: READ <= 8'Hf1;
      32'H229: READ <= 8'Hf2;
      32'H230: READ <= 8'Hf2;
      32'H231: READ <= 8'Hf2;
      32'H232: READ <= 8'Hf2;
      32'H233: READ <= 8'Hf2;
      32'H234: READ <= 8'Hf2;
      32'H235: READ <= 8'Hf1;
      32'H236: READ <= 8'Hef;
      32'H237: READ <= 8'Hee;
      32'H238: READ <= 8'Hed;
      32'H239: READ <= 8'Hec;
      32'H240: READ <= 8'Hea;
      32'H241: READ <= 8'Heb;
      32'H242: READ <= 8'Hea;
      32'H243: READ <= 8'He6;
      32'H244: READ <= 8'He1;
      32'H245: READ <= 8'Hdd;
      32'H246: READ <= 8'Hda;
      32'H247: READ <= 8'Hd5;
      32'H248: READ <= 8'Hd1;
      32'H249: READ <= 8'Hcc;
      32'H250: READ <= 8'Hc6;
      32'H251: READ <= 8'Hbe;
      32'H252: READ <= 8'Hb6;
      32'H253: READ <= 8'Had;
      32'H254: READ <= 8'Ha7;
      32'H255: READ <= 8'Ha1;
      32'H256: READ <= 8'H9e;
      32'H257: READ <= 8'H9c;
      32'H258: READ <= 8'H9a;
      32'H259: READ <= 8'H9a;
      32'H260: READ <= 8'H98;
      32'H261: READ <= 8'H98;
      32'H262: READ <= 8'H98;
      32'H263: READ <= 8'H98;
      32'H264: READ <= 8'H99;
      32'H265: READ <= 8'H99;
      32'H266: READ <= 8'H99;
      32'H267: READ <= 8'H9a;
      32'H268: READ <= 8'H9a;
      32'H269: READ <= 8'H9b;
      32'H270: READ <= 8'H9b;
      32'H271: READ <= 8'H9b;
      32'H272: READ <= 8'H9a;
      32'H273: READ <= 8'H9b;
      32'H274: READ <= 8'H9b;
      32'H275: READ <= 8'H9c;
      32'H276: READ <= 8'H9d;
      32'H277: READ <= 8'H9d;
      32'H278: READ <= 8'H9e;
      32'H279: READ <= 8'H9e;
      32'H280: READ <= 8'H9f;
      32'H281: READ <= 8'H9f;
      32'H282: READ <= 8'Ha0;
      32'H283: READ <= 8'Ha1;
      32'H284: READ <= 8'Ha2;
      32'H285: READ <= 8'Ha1;
      32'H286: READ <= 8'Ha1;
      32'H287: READ <= 8'Ha2;
      32'H288: READ <= 8'Ha1;
      32'H289: READ <= 8'Ha2;
      32'H290: READ <= 8'Ha2;
      32'H291: READ <= 8'Ha1;
      32'H292: READ <= 8'Ha2;
      32'H293: READ <= 8'Ha3;
      32'H294: READ <= 8'Ha3;
      32'H295: READ <= 8'Ha3;
      32'H296: READ <= 8'Ha4;
      32'H297: READ <= 8'Ha5;
      32'H298: READ <= 8'Ha5;
      32'H299: READ <= 8'Ha6;
      32'H300: READ <= 8'Haf;
      32'H301: READ <= 8'Hb3;
      32'H302: READ <= 8'Hb5;
      32'H303: READ <= 8'Hb6;
      32'H304: READ <= 8'Hb9;
      32'H305: READ <= 8'Hbb;
      32'H306: READ <= 8'Hbf;
      32'H307: READ <= 8'Hc3;
      32'H308: READ <= 8'Hc6;
      32'H309: READ <= 8'Hca;
      32'H310: READ <= 8'Hcd;
      32'H311: READ <= 8'Hd1;
      32'H312: READ <= 8'Hd3;
      32'H313: READ <= 8'Hd6;
      32'H314: READ <= 8'Hda;
      32'H315: READ <= 8'Hdc;
      32'H316: READ <= 8'Hdf;
      32'H317: READ <= 8'He2;
      32'H318: READ <= 8'He5;
      32'H319: READ <= 8'He7;
      32'H320: READ <= 8'He8;
      32'H321: READ <= 8'Hea;
      32'H322: READ <= 8'Heb;
      32'H323: READ <= 8'Heb;
      32'H324: READ <= 8'Hed;
      32'H325: READ <= 8'Hee;
      32'H326: READ <= 8'Hee;
      32'H327: READ <= 8'Hf0;
      32'H328: READ <= 8'Hf1;
      32'H329: READ <= 8'Hf2;
      32'H330: READ <= 8'Hf2;
      32'H331: READ <= 8'Hf3;
      32'H332: READ <= 8'Hf3;
      32'H333: READ <= 8'Hf2;
      32'H334: READ <= 8'Hf2;
      32'H335: READ <= 8'Hf1;
      32'H336: READ <= 8'Hef;
      32'H337: READ <= 8'Hee;
      32'H338: READ <= 8'Hed;
      32'H339: READ <= 8'Hed;
      32'H340: READ <= 8'Hed;
      32'H341: READ <= 8'Hee;
      32'H342: READ <= 8'Hee;
      32'H343: READ <= 8'Hec;
      32'H344: READ <= 8'He3;
      32'H345: READ <= 8'Hde;
      32'H346: READ <= 8'Hdb;
      32'H347: READ <= 8'Hd7;
      32'H348: READ <= 8'Hd1;
      32'H349: READ <= 8'Hcd;
      32'H350: READ <= 8'Hc7;
      32'H351: READ <= 8'Hc0;
      32'H352: READ <= 8'Hb7;
      32'H353: READ <= 8'Haf;
      32'H354: READ <= 8'Ha7;
      32'H355: READ <= 8'Ha2;
      32'H356: READ <= 8'H9e;
      32'H357: READ <= 8'H9b;
      32'H358: READ <= 8'H9a;
      32'H359: READ <= 8'H99;
      32'H360: READ <= 8'H97;
      32'H361: READ <= 8'H96;
      32'H362: READ <= 8'H97;
      32'H363: READ <= 8'H97;
      32'H364: READ <= 8'H97;
      32'H365: READ <= 8'H98;
      32'H366: READ <= 8'H98;
      32'H367: READ <= 8'H99;
      32'H368: READ <= 8'H99;
      32'H369: READ <= 8'H9a;
      32'H370: READ <= 8'H9a;
      32'H371: READ <= 8'H9a;
      32'H372: READ <= 8'H99;
      32'H373: READ <= 8'H9a;
      32'H374: READ <= 8'H9a;
      32'H375: READ <= 8'H9b;
      32'H376: READ <= 8'H9b;
      32'H377: READ <= 8'H9c;
      32'H378: READ <= 8'H9d;
      32'H379: READ <= 8'H9e;
      32'H380: READ <= 8'H9e;
      32'H381: READ <= 8'H9f;
      32'H382: READ <= 8'H9f;
      32'H383: READ <= 8'Ha0;
      32'H384: READ <= 8'Ha0;
      32'H385: READ <= 8'Ha0;
      32'H386: READ <= 8'Ha0;
      32'H387: READ <= 8'Ha1;
      32'H388: READ <= 8'Ha1;
      32'H389: READ <= 8'Ha1;
      32'H390: READ <= 8'Ha1;
      32'H391: READ <= 8'Ha1;
      32'H392: READ <= 8'Ha1;
      32'H393: READ <= 8'Ha1;
      32'H394: READ <= 8'Ha1;
      32'H395: READ <= 8'Ha2;
      32'H396: READ <= 8'Ha3;
      32'H397: READ <= 8'Ha4;
      32'H398: READ <= 8'Ha4;
      32'H399: READ <= 8'Ha5;
      32'H400: READ <= 8'Had;
      32'H401: READ <= 8'Hb1;
      32'H402: READ <= 8'Hb3;
      32'H403: READ <= 8'Hb4;
      32'H404: READ <= 8'Hb6;
      32'H405: READ <= 8'Hba;
      32'H406: READ <= 8'Hbe;
      32'H407: READ <= 8'Hc1;
      32'H408: READ <= 8'Hc4;
      32'H409: READ <= 8'Hc8;
      32'H410: READ <= 8'Hcc;
      32'H411: READ <= 8'Hd0;
      32'H412: READ <= 8'Hd2;
      32'H413: READ <= 8'Hd5;
      32'H414: READ <= 8'Hd8;
      32'H415: READ <= 8'Hdc;
      32'H416: READ <= 8'Hdf;
      32'H417: READ <= 8'He1;
      32'H418: READ <= 8'He4;
      32'H419: READ <= 8'He7;
      32'H420: READ <= 8'He8;
      32'H421: READ <= 8'He9;
      32'H422: READ <= 8'Heb;
      32'H423: READ <= 8'Hec;
      32'H424: READ <= 8'Hed;
      32'H425: READ <= 8'Hee;
      32'H426: READ <= 8'Hef;
      32'H427: READ <= 8'Hf0;
      32'H428: READ <= 8'Hf1;
      32'H429: READ <= 8'Hf2;
      32'H430: READ <= 8'Hf2;
      32'H431: READ <= 8'Hf2;
      32'H432: READ <= 8'Hf3;
      32'H433: READ <= 8'Hf2;
      32'H434: READ <= 8'Hf2;
      32'H435: READ <= 8'Hf1;
      32'H436: READ <= 8'Hf0;
      32'H437: READ <= 8'Hf0;
      32'H438: READ <= 8'Hf0;
      32'H439: READ <= 8'Hef;
      32'H440: READ <= 8'Heb;
      32'H441: READ <= 8'He4;
      32'H442: READ <= 8'Hdc;
      32'H443: READ <= 8'Hdf;
      32'H444: READ <= 8'He2;
      32'H445: READ <= 8'He4;
      32'H446: READ <= 8'He1;
      32'H447: READ <= 8'Hde;
      32'H448: READ <= 8'Hda;
      32'H449: READ <= 8'Hd1;
      32'H450: READ <= 8'Hcc;
      32'H451: READ <= 8'Hc2;
      32'H452: READ <= 8'Hb9;
      32'H453: READ <= 8'Haf;
      32'H454: READ <= 8'Ha8;
      32'H455: READ <= 8'Ha2;
      32'H456: READ <= 8'H9e;
      32'H457: READ <= 8'H9a;
      32'H458: READ <= 8'H99;
      32'H459: READ <= 8'H98;
      32'H460: READ <= 8'H98;
      32'H461: READ <= 8'H96;
      32'H462: READ <= 8'H96;
      32'H463: READ <= 8'H96;
      32'H464: READ <= 8'H95;
      32'H465: READ <= 8'H96;
      32'H466: READ <= 8'H97;
      32'H467: READ <= 8'H97;
      32'H468: READ <= 8'H98;
      32'H469: READ <= 8'H99;
      32'H470: READ <= 8'H99;
      32'H471: READ <= 8'H99;
      32'H472: READ <= 8'H99;
      32'H473: READ <= 8'H99;
      32'H474: READ <= 8'H99;
      32'H475: READ <= 8'H9a;
      32'H476: READ <= 8'H99;
      32'H477: READ <= 8'H9b;
      32'H478: READ <= 8'H9c;
      32'H479: READ <= 8'H9c;
      32'H480: READ <= 8'H9d;
      32'H481: READ <= 8'H9e;
      32'H482: READ <= 8'H9d;
      32'H483: READ <= 8'H9e;
      32'H484: READ <= 8'H9e;
      32'H485: READ <= 8'H9f;
      32'H486: READ <= 8'H9f;
      32'H487: READ <= 8'H9f;
      32'H488: READ <= 8'Ha0;
      32'H489: READ <= 8'Ha0;
      32'H490: READ <= 8'Ha0;
      32'H491: READ <= 8'Ha1;
      32'H492: READ <= 8'Ha0;
      32'H493: READ <= 8'Ha0;
      32'H494: READ <= 8'Ha1;
      32'H495: READ <= 8'Ha2;
      32'H496: READ <= 8'Ha2;
      32'H497: READ <= 8'Ha2;
      32'H498: READ <= 8'Ha3;
      32'H499: READ <= 8'Ha4;
      32'H500: READ <= 8'Hab;
      32'H501: READ <= 8'Haf;
      32'H502: READ <= 8'Hb1;
      32'H503: READ <= 8'Hb3;
      32'H504: READ <= 8'Hb5;
      32'H505: READ <= 8'Hb8;
      32'H506: READ <= 8'Hbb;
      32'H507: READ <= 8'Hbf;
      32'H508: READ <= 8'Hc2;
      32'H509: READ <= 8'Hc6;
      32'H510: READ <= 8'Hcb;
      32'H511: READ <= 8'Hce;
      32'H512: READ <= 8'Hd2;
      32'H513: READ <= 8'Hd4;
      32'H514: READ <= 8'Hd7;
      32'H515: READ <= 8'Hdb;
      32'H516: READ <= 8'Hde;
      32'H517: READ <= 8'He1;
      32'H518: READ <= 8'He4;
      32'H519: READ <= 8'He6;
      32'H520: READ <= 8'He8;
      32'H521: READ <= 8'He9;
      32'H522: READ <= 8'Heb;
      32'H523: READ <= 8'Hec;
      32'H524: READ <= 8'Hed;
      32'H525: READ <= 8'Hee;
      32'H526: READ <= 8'Hef;
      32'H527: READ <= 8'Hf1;
      32'H528: READ <= 8'Hf1;
      32'H529: READ <= 8'Hf2;
      32'H530: READ <= 8'Hf3;
      32'H531: READ <= 8'Hf3;
      32'H532: READ <= 8'Hf3;
      32'H533: READ <= 8'Hf2;
      32'H534: READ <= 8'Hf3;
      32'H535: READ <= 8'Hf1;
      32'H536: READ <= 8'Hf4;
      32'H537: READ <= 8'Hef;
      32'H538: READ <= 8'Hd5;
      32'H539: READ <= 8'Hca;
      32'H540: READ <= 8'Hc2;
      32'H541: READ <= 8'Hc2;
      32'H542: READ <= 8'Hbd;
      32'H543: READ <= 8'Hb6;
      32'H544: READ <= 8'Hbc;
      32'H545: READ <= 8'Hc6;
      32'H546: READ <= 8'Hcc;
      32'H547: READ <= 8'Hbc;
      32'H548: READ <= 8'Hc1;
      32'H549: READ <= 8'Hc8;
      32'H550: READ <= 8'Hba;
      32'H551: READ <= 8'Hc2;
      32'H552: READ <= 8'Hb8;
      32'H553: READ <= 8'Hb1;
      32'H554: READ <= 8'Ha9;
      32'H555: READ <= 8'Ha2;
      32'H556: READ <= 8'H9d;
      32'H557: READ <= 8'H9a;
      32'H558: READ <= 8'H98;
      32'H559: READ <= 8'H97;
      32'H560: READ <= 8'H97;
      32'H561: READ <= 8'H95;
      32'H562: READ <= 8'H95;
      32'H563: READ <= 8'H95;
      32'H564: READ <= 8'H95;
      32'H565: READ <= 8'H96;
      32'H566: READ <= 8'H96;
      32'H567: READ <= 8'H96;
      32'H568: READ <= 8'H97;
      32'H569: READ <= 8'H98;
      32'H570: READ <= 8'H97;
      32'H571: READ <= 8'H97;
      32'H572: READ <= 8'H97;
      32'H573: READ <= 8'H98;
      32'H574: READ <= 8'H98;
      32'H575: READ <= 8'H99;
      32'H576: READ <= 8'H99;
      32'H577: READ <= 8'H9a;
      32'H578: READ <= 8'H9b;
      32'H579: READ <= 8'H9c;
      32'H580: READ <= 8'H9c;
      32'H581: READ <= 8'H9d;
      32'H582: READ <= 8'H9d;
      32'H583: READ <= 8'H9d;
      32'H584: READ <= 8'H9d;
      32'H585: READ <= 8'H9e;
      32'H586: READ <= 8'H9e;
      32'H587: READ <= 8'H9e;
      32'H588: READ <= 8'H9f;
      32'H589: READ <= 8'H9f;
      32'H590: READ <= 8'H9f;
      32'H591: READ <= 8'Ha0;
      32'H592: READ <= 8'Ha0;
      32'H593: READ <= 8'Ha0;
      32'H594: READ <= 8'Ha0;
      32'H595: READ <= 8'Ha0;
      32'H596: READ <= 8'Ha1;
      32'H597: READ <= 8'Ha2;
      32'H598: READ <= 8'Ha2;
      32'H599: READ <= 8'Ha2;
      32'H600: READ <= 8'Ha9;
      32'H601: READ <= 8'Hac;
      32'H602: READ <= 8'Haf;
      32'H603: READ <= 8'Hb2;
      32'H604: READ <= 8'Hb4;
      32'H605: READ <= 8'Hb7;
      32'H606: READ <= 8'Hba;
      32'H607: READ <= 8'Hbd;
      32'H608: READ <= 8'Hc1;
      32'H609: READ <= 8'Hc4;
      32'H610: READ <= 8'Hc9;
      32'H611: READ <= 8'Hcd;
      32'H612: READ <= 8'Hd1;
      32'H613: READ <= 8'Hd3;
      32'H614: READ <= 8'Hd6;
      32'H615: READ <= 8'Hd9;
      32'H616: READ <= 8'Hdd;
      32'H617: READ <= 8'He0;
      32'H618: READ <= 8'He3;
      32'H619: READ <= 8'He5;
      32'H620: READ <= 8'He7;
      32'H621: READ <= 8'He9;
      32'H622: READ <= 8'Heb;
      32'H623: READ <= 8'Hec;
      32'H624: READ <= 8'Hed;
      32'H625: READ <= 8'Hee;
      32'H626: READ <= 8'Hef;
      32'H627: READ <= 8'Hf0;
      32'H628: READ <= 8'Hf1;
      32'H629: READ <= 8'Hf2;
      32'H630: READ <= 8'Hf3;
      32'H631: READ <= 8'Hf3;
      32'H632: READ <= 8'Hf3;
      32'H633: READ <= 8'Hf3;
      32'H634: READ <= 8'Hf1;
      32'H635: READ <= 8'Hf8;
      32'H636: READ <= 8'He5;
      32'H637: READ <= 8'Hbb;
      32'H638: READ <= 8'H9e;
      32'H639: READ <= 8'Haa;
      32'H640: READ <= 8'Hb3;
      32'H641: READ <= 8'Ha8;
      32'H642: READ <= 8'Had;
      32'H643: READ <= 8'Hac;
      32'H644: READ <= 8'H9e;
      32'H645: READ <= 8'Ha3;
      32'H646: READ <= 8'H9b;
      32'H647: READ <= 8'H9e;
      32'H648: READ <= 8'H93;
      32'H649: READ <= 8'Ha7;
      32'H650: READ <= 8'Ha1;
      32'H651: READ <= 8'H9e;
      32'H652: READ <= 8'Hac;
      32'H653: READ <= 8'Hb6;
      32'H654: READ <= 8'Hac;
      32'H655: READ <= 8'Ha2;
      32'H656: READ <= 8'H9d;
      32'H657: READ <= 8'H99;
      32'H658: READ <= 8'H98;
      32'H659: READ <= 8'H96;
      32'H660: READ <= 8'H96;
      32'H661: READ <= 8'H95;
      32'H662: READ <= 8'H94;
      32'H663: READ <= 8'H94;
      32'H664: READ <= 8'H93;
      32'H665: READ <= 8'H94;
      32'H666: READ <= 8'H95;
      32'H667: READ <= 8'H95;
      32'H668: READ <= 8'H96;
      32'H669: READ <= 8'H96;
      32'H670: READ <= 8'H96;
      32'H671: READ <= 8'H96;
      32'H672: READ <= 8'H96;
      32'H673: READ <= 8'H97;
      32'H674: READ <= 8'H97;
      32'H675: READ <= 8'H97;
      32'H676: READ <= 8'H99;
      32'H677: READ <= 8'H99;
      32'H678: READ <= 8'H9a;
      32'H679: READ <= 8'H9b;
      32'H680: READ <= 8'H9b;
      32'H681: READ <= 8'H9b;
      32'H682: READ <= 8'H9c;
      32'H683: READ <= 8'H9c;
      32'H684: READ <= 8'H9c;
      32'H685: READ <= 8'H9e;
      32'H686: READ <= 8'H9e;
      32'H687: READ <= 8'H9e;
      32'H688: READ <= 8'H9e;
      32'H689: READ <= 8'H9e;
      32'H690: READ <= 8'H9f;
      32'H691: READ <= 8'H9f;
      32'H692: READ <= 8'H9e;
      32'H693: READ <= 8'H9e;
      32'H694: READ <= 8'H9f;
      32'H695: READ <= 8'H9f;
      32'H696: READ <= 8'Ha0;
      32'H697: READ <= 8'Ha1;
      32'H698: READ <= 8'Ha1;
      32'H699: READ <= 8'Ha1;
      32'H700: READ <= 8'Ha7;
      32'H701: READ <= 8'Ha9;
      32'H702: READ <= 8'Had;
      32'H703: READ <= 8'Hb0;
      32'H704: READ <= 8'Hb2;
      32'H705: READ <= 8'Hb6;
      32'H706: READ <= 8'Hb8;
      32'H707: READ <= 8'Hbc;
      32'H708: READ <= 8'Hc0;
      32'H709: READ <= 8'Hc2;
      32'H710: READ <= 8'Hc7;
      32'H711: READ <= 8'Hcc;
      32'H712: READ <= 8'Hd0;
      32'H713: READ <= 8'Hd2;
      32'H714: READ <= 8'Hd5;
      32'H715: READ <= 8'Hd8;
      32'H716: READ <= 8'Hdc;
      32'H717: READ <= 8'Hdf;
      32'H718: READ <= 8'He2;
      32'H719: READ <= 8'He5;
      32'H720: READ <= 8'He7;
      32'H721: READ <= 8'He8;
      32'H722: READ <= 8'Hea;
      32'H723: READ <= 8'Heb;
      32'H724: READ <= 8'Hed;
      32'H725: READ <= 8'Hee;
      32'H726: READ <= 8'Hef;
      32'H727: READ <= 8'Hf0;
      32'H728: READ <= 8'Hf1;
      32'H729: READ <= 8'Hf2;
      32'H730: READ <= 8'Hf2;
      32'H731: READ <= 8'Hf3;
      32'H732: READ <= 8'Hf3;
      32'H733: READ <= 8'Hf5;
      32'H734: READ <= 8'Hf7;
      32'H735: READ <= 8'Hc8;
      32'H736: READ <= 8'Ha8;
      32'H737: READ <= 8'Haa;
      32'H738: READ <= 8'Ha1;
      32'H739: READ <= 8'H88;
      32'H740: READ <= 8'Hae;
      32'H741: READ <= 8'Ha6;
      32'H742: READ <= 8'Hac;
      32'H743: READ <= 8'Ha3;
      32'H744: READ <= 8'H99;
      32'H745: READ <= 8'H93;
      32'H746: READ <= 8'H91;
      32'H747: READ <= 8'H93;
      32'H748: READ <= 8'H82;
      32'H749: READ <= 8'H92;
      32'H750: READ <= 8'H85;
      32'H751: READ <= 8'H77;
      32'H752: READ <= 8'H83;
      32'H753: READ <= 8'H9b;
      32'H754: READ <= 8'Hb2;
      32'H755: READ <= 8'Ha7;
      32'H756: READ <= 8'H9d;
      32'H757: READ <= 8'H9a;
      32'H758: READ <= 8'H97;
      32'H759: READ <= 8'H96;
      32'H760: READ <= 8'H95;
      32'H761: READ <= 8'H94;
      32'H762: READ <= 8'H93;
      32'H763: READ <= 8'H92;
      32'H764: READ <= 8'H93;
      32'H765: READ <= 8'H93;
      32'H766: READ <= 8'H94;
      32'H767: READ <= 8'H94;
      32'H768: READ <= 8'H94;
      32'H769: READ <= 8'H95;
      32'H770: READ <= 8'H95;
      32'H771: READ <= 8'H95;
      32'H772: READ <= 8'H95;
      32'H773: READ <= 8'H96;
      32'H774: READ <= 8'H97;
      32'H775: READ <= 8'H97;
      32'H776: READ <= 8'H96;
      32'H777: READ <= 8'H98;
      32'H778: READ <= 8'H99;
      32'H779: READ <= 8'H9a;
      32'H780: READ <= 8'H9a;
      32'H781: READ <= 8'H9b;
      32'H782: READ <= 8'H9b;
      32'H783: READ <= 8'H9c;
      32'H784: READ <= 8'H9d;
      32'H785: READ <= 8'H9d;
      32'H786: READ <= 8'H9d;
      32'H787: READ <= 8'H9d;
      32'H788: READ <= 8'H9d;
      32'H789: READ <= 8'H9d;
      32'H790: READ <= 8'H9e;
      32'H791: READ <= 8'H9e;
      32'H792: READ <= 8'H9e;
      32'H793: READ <= 8'H9e;
      32'H794: READ <= 8'H9d;
      32'H795: READ <= 8'H9e;
      32'H796: READ <= 8'H9e;
      32'H797: READ <= 8'H9f;
      32'H798: READ <= 8'Ha0;
      32'H799: READ <= 8'Ha0;
      32'H800: READ <= 8'Ha5;
      32'H801: READ <= 8'Ha7;
      32'H802: READ <= 8'Hab;
      32'H803: READ <= 8'Haf;
      32'H804: READ <= 8'Hb1;
      32'H805: READ <= 8'Hb5;
      32'H806: READ <= 8'Hb7;
      32'H807: READ <= 8'Hbb;
      32'H808: READ <= 8'Hbd;
      32'H809: READ <= 8'Hc1;
      32'H810: READ <= 8'Hc5;
      32'H811: READ <= 8'Hca;
      32'H812: READ <= 8'Hcc;
      32'H813: READ <= 8'Hd0;
      32'H814: READ <= 8'Hd4;
      32'H815: READ <= 8'Hd7;
      32'H816: READ <= 8'Hdb;
      32'H817: READ <= 8'Hde;
      32'H818: READ <= 8'He1;
      32'H819: READ <= 8'He4;
      32'H820: READ <= 8'He6;
      32'H821: READ <= 8'He9;
      32'H822: READ <= 8'Hea;
      32'H823: READ <= 8'Heb;
      32'H824: READ <= 8'Hed;
      32'H825: READ <= 8'Hee;
      32'H826: READ <= 8'Hef;
      32'H827: READ <= 8'Hf0;
      32'H828: READ <= 8'Hf2;
      32'H829: READ <= 8'Hf2;
      32'H830: READ <= 8'Hf3;
      32'H831: READ <= 8'Hf3;
      32'H832: READ <= 8'Hee;
      32'H833: READ <= 8'Hc2;
      32'H834: READ <= 8'H9c;
      32'H835: READ <= 8'H60;
      32'H836: READ <= 8'H62;
      32'H837: READ <= 8'H64;
      32'H838: READ <= 8'H7a;
      32'H839: READ <= 8'H83;
      32'H840: READ <= 8'H99;
      32'H841: READ <= 8'H97;
      32'H842: READ <= 8'H98;
      32'H843: READ <= 8'Haf;
      32'H844: READ <= 8'H96;
      32'H845: READ <= 8'H92;
      32'H846: READ <= 8'H9a;
      32'H847: READ <= 8'H9e;
      32'H848: READ <= 8'H81;
      32'H849: READ <= 8'H8b;
      32'H850: READ <= 8'H79;
      32'H851: READ <= 8'H8b;
      32'H852: READ <= 8'H82;
      32'H853: READ <= 8'H9a;
      32'H854: READ <= 8'H9e;
      32'H855: READ <= 8'Ha9;
      32'H856: READ <= 8'H9e;
      32'H857: READ <= 8'H99;
      32'H858: READ <= 8'H98;
      32'H859: READ <= 8'H96;
      32'H860: READ <= 8'H95;
      32'H861: READ <= 8'H93;
      32'H862: READ <= 8'H91;
      32'H863: READ <= 8'H91;
      32'H864: READ <= 8'H92;
      32'H865: READ <= 8'H92;
      32'H866: READ <= 8'H92;
      32'H867: READ <= 8'H93;
      32'H868: READ <= 8'H92;
      32'H869: READ <= 8'H93;
      32'H870: READ <= 8'H93;
      32'H871: READ <= 8'H94;
      32'H872: READ <= 8'H94;
      32'H873: READ <= 8'H95;
      32'H874: READ <= 8'H94;
      32'H875: READ <= 8'H96;
      32'H876: READ <= 8'H95;
      32'H877: READ <= 8'H96;
      32'H878: READ <= 8'H98;
      32'H879: READ <= 8'H99;
      32'H880: READ <= 8'H99;
      32'H881: READ <= 8'H99;
      32'H882: READ <= 8'H9a;
      32'H883: READ <= 8'H9b;
      32'H884: READ <= 8'H9b;
      32'H885: READ <= 8'H9c;
      32'H886: READ <= 8'H9d;
      32'H887: READ <= 8'H9c;
      32'H888: READ <= 8'H9c;
      32'H889: READ <= 8'H9c;
      32'H890: READ <= 8'H9c;
      32'H891: READ <= 8'H9d;
      32'H892: READ <= 8'H9d;
      32'H893: READ <= 8'H9c;
      32'H894: READ <= 8'H9d;
      32'H895: READ <= 8'H9c;
      32'H896: READ <= 8'H9d;
      32'H897: READ <= 8'H9e;
      32'H898: READ <= 8'H9e;
      32'H899: READ <= 8'H9f;
      32'H900: READ <= 8'Ha4;
      32'H901: READ <= 8'Ha7;
      32'H902: READ <= 8'Ha9;
      32'H903: READ <= 8'Had;
      32'H904: READ <= 8'Hb0;
      32'H905: READ <= 8'Hb3;
      32'H906: READ <= 8'Hb5;
      32'H907: READ <= 8'Hb9;
      32'H908: READ <= 8'Hbb;
      32'H909: READ <= 8'Hbf;
      32'H910: READ <= 8'Hc3;
      32'H911: READ <= 8'Hc7;
      32'H912: READ <= 8'Hcb;
      32'H913: READ <= 8'Hcf;
      32'H914: READ <= 8'Hd2;
      32'H915: READ <= 8'Hd6;
      32'H916: READ <= 8'Hd9;
      32'H917: READ <= 8'Hdd;
      32'H918: READ <= 8'He0;
      32'H919: READ <= 8'He4;
      32'H920: READ <= 8'He6;
      32'H921: READ <= 8'He7;
      32'H922: READ <= 8'Hea;
      32'H923: READ <= 8'Hec;
      32'H924: READ <= 8'Hed;
      32'H925: READ <= 8'Hed;
      32'H926: READ <= 8'Hf0;
      32'H927: READ <= 8'Hf1;
      32'H928: READ <= 8'Hf1;
      32'H929: READ <= 8'Hf3;
      32'H930: READ <= 8'Hf1;
      32'H931: READ <= 8'Hcb;
      32'H932: READ <= 8'Ha5;
      32'H933: READ <= 8'H88;
      32'H934: READ <= 8'H75;
      32'H935: READ <= 8'H81;
      32'H936: READ <= 8'H8c;
      32'H937: READ <= 8'H4a;
      32'H938: READ <= 8'H5f;
      32'H939: READ <= 8'Ha1;
      32'H940: READ <= 8'Ha6;
      32'H941: READ <= 8'H90;
      32'H942: READ <= 8'H93;
      32'H943: READ <= 8'H96;
      32'H944: READ <= 8'H93;
      32'H945: READ <= 8'H96;
      32'H946: READ <= 8'H9e;
      32'H947: READ <= 8'Hb1;
      32'H948: READ <= 8'H67;
      32'H949: READ <= 8'H7f;
      32'H950: READ <= 8'Hb0;
      32'H951: READ <= 8'Hc2;
      32'H952: READ <= 8'Hd8;
      32'H953: READ <= 8'Hdb;
      32'H954: READ <= 8'Hbd;
      32'H955: READ <= 8'Ha9;
      32'H956: READ <= 8'Hac;
      32'H957: READ <= 8'H9f;
      32'H958: READ <= 8'H99;
      32'H959: READ <= 8'H96;
      32'H960: READ <= 8'H95;
      32'H961: READ <= 8'H93;
      32'H962: READ <= 8'H91;
      32'H963: READ <= 8'H90;
      32'H964: READ <= 8'H90;
      32'H965: READ <= 8'H90;
      32'H966: READ <= 8'H91;
      32'H967: READ <= 8'H92;
      32'H968: READ <= 8'H92;
      32'H969: READ <= 8'H92;
      32'H970: READ <= 8'H92;
      32'H971: READ <= 8'H92;
      32'H972: READ <= 8'H92;
      32'H973: READ <= 8'H93;
      32'H974: READ <= 8'H93;
      32'H975: READ <= 8'H95;
      32'H976: READ <= 8'H95;
      32'H977: READ <= 8'H95;
      32'H978: READ <= 8'H97;
      32'H979: READ <= 8'H99;
      32'H980: READ <= 8'H98;
      32'H981: READ <= 8'H99;
      32'H982: READ <= 8'H9a;
      32'H983: READ <= 8'H9a;
      32'H984: READ <= 8'H9a;
      32'H985: READ <= 8'H9a;
      32'H986: READ <= 8'H9b;
      32'H987: READ <= 8'H9b;
      32'H988: READ <= 8'H9c;
      32'H989: READ <= 8'H9c;
      32'H990: READ <= 8'H9b;
      32'H991: READ <= 8'H9c;
      32'H992: READ <= 8'H9b;
      32'H993: READ <= 8'H9c;
      32'H994: READ <= 8'H9c;
      32'H995: READ <= 8'H9c;
      32'H996: READ <= 8'H9d;
      32'H997: READ <= 8'H9d;
      32'H998: READ <= 8'H9d;
      32'H999: READ <= 8'H9e;
      32'H1000: READ <= 8'Ha3;
      32'H1001: READ <= 8'Ha5;
      32'H1002: READ <= 8'Ha8;
      32'H1003: READ <= 8'Hab;
      32'H1004: READ <= 8'Hae;
      32'H1005: READ <= 8'Hb1;
      32'H1006: READ <= 8'Hb5;
      32'H1007: READ <= 8'Hb6;
      32'H1008: READ <= 8'Hba;
      32'H1009: READ <= 8'Hbd;
      32'H1010: READ <= 8'Hc0;
      32'H1011: READ <= 8'Hc5;
      32'H1012: READ <= 8'Hc9;
      32'H1013: READ <= 8'Hcd;
      32'H1014: READ <= 8'Hcf;
      32'H1015: READ <= 8'Hd3;
      32'H1016: READ <= 8'Hd7;
      32'H1017: READ <= 8'Hdb;
      32'H1018: READ <= 8'Hdf;
      32'H1019: READ <= 8'He2;
      32'H1020: READ <= 8'He4;
      32'H1021: READ <= 8'He7;
      32'H1022: READ <= 8'He9;
      32'H1023: READ <= 8'Heb;
      32'H1024: READ <= 8'Hec;
      32'H1025: READ <= 8'Hed;
      32'H1026: READ <= 8'Hef;
      32'H1027: READ <= 8'Hf2;
      32'H1028: READ <= 8'Hf2;
      32'H1029: READ <= 8'He6;
      32'H1030: READ <= 8'Haf;
      32'H1031: READ <= 8'H92;
      32'H1032: READ <= 8'H7f;
      32'H1033: READ <= 8'H8c;
      32'H1034: READ <= 8'H90;
      32'H1035: READ <= 8'H8a;
      32'H1036: READ <= 8'H8b;
      32'H1037: READ <= 8'H85;
      32'H1038: READ <= 8'H33;
      32'H1039: READ <= 8'H76;
      32'H1040: READ <= 8'H8e;
      32'H1041: READ <= 8'H96;
      32'H1042: READ <= 8'H81;
      32'H1043: READ <= 8'H88;
      32'H1044: READ <= 8'H97;
      32'H1045: READ <= 8'Ha3;
      32'H1046: READ <= 8'Hae;
      32'H1047: READ <= 8'H7a;
      32'H1048: READ <= 8'H9f;
      32'H1049: READ <= 8'Hc9;
      32'H1050: READ <= 8'Hd5;
      32'H1051: READ <= 8'Hde;
      32'H1052: READ <= 8'Hde;
      32'H1053: READ <= 8'Hda;
      32'H1054: READ <= 8'Hc1;
      32'H1055: READ <= 8'Haa;
      32'H1056: READ <= 8'Had;
      32'H1057: READ <= 8'H9a;
      32'H1058: READ <= 8'Ha0;
      32'H1059: READ <= 8'H9b;
      32'H1060: READ <= 8'H96;
      32'H1061: READ <= 8'H93;
      32'H1062: READ <= 8'H91;
      32'H1063: READ <= 8'H8f;
      32'H1064: READ <= 8'H8f;
      32'H1065: READ <= 8'H8e;
      32'H1066: READ <= 8'H90;
      32'H1067: READ <= 8'H90;
      32'H1068: READ <= 8'H91;
      32'H1069: READ <= 8'H91;
      32'H1070: READ <= 8'H90;
      32'H1071: READ <= 8'H92;
      32'H1072: READ <= 8'H92;
      32'H1073: READ <= 8'H91;
      32'H1074: READ <= 8'H93;
      32'H1075: READ <= 8'H93;
      32'H1076: READ <= 8'H94;
      32'H1077: READ <= 8'H96;
      32'H1078: READ <= 8'H97;
      32'H1079: READ <= 8'H97;
      32'H1080: READ <= 8'H98;
      32'H1081: READ <= 8'H98;
      32'H1082: READ <= 8'H98;
      32'H1083: READ <= 8'H99;
      32'H1084: READ <= 8'H99;
      32'H1085: READ <= 8'H99;
      32'H1086: READ <= 8'H99;
      32'H1087: READ <= 8'H9b;
      32'H1088: READ <= 8'H9b;
      32'H1089: READ <= 8'H9a;
      32'H1090: READ <= 8'H9a;
      32'H1091: READ <= 8'H9b;
      32'H1092: READ <= 8'H9b;
      32'H1093: READ <= 8'H9a;
      32'H1094: READ <= 8'H9a;
      32'H1095: READ <= 8'H9b;
      32'H1096: READ <= 8'H9b;
      32'H1097: READ <= 8'H9c;
      32'H1098: READ <= 8'H9c;
      32'H1099: READ <= 8'H9d;
      32'H1100: READ <= 8'Ha1;
      32'H1101: READ <= 8'Ha3;
      32'H1102: READ <= 8'Ha6;
      32'H1103: READ <= 8'Ha9;
      32'H1104: READ <= 8'Had;
      32'H1105: READ <= 8'Hb0;
      32'H1106: READ <= 8'Hb2;
      32'H1107: READ <= 8'Hb4;
      32'H1108: READ <= 8'Hb8;
      32'H1109: READ <= 8'Hbc;
      32'H1110: READ <= 8'Hbe;
      32'H1111: READ <= 8'Hc2;
      32'H1112: READ <= 8'Hc7;
      32'H1113: READ <= 8'Hcb;
      32'H1114: READ <= 8'Hcd;
      32'H1115: READ <= 8'Hd1;
      32'H1116: READ <= 8'Hd6;
      32'H1117: READ <= 8'Hd9;
      32'H1118: READ <= 8'Hdc;
      32'H1119: READ <= 8'He0;
      32'H1120: READ <= 8'He4;
      32'H1121: READ <= 8'He6;
      32'H1122: READ <= 8'He9;
      32'H1123: READ <= 8'Heb;
      32'H1124: READ <= 8'Hec;
      32'H1125: READ <= 8'Hed;
      32'H1126: READ <= 8'Hef;
      32'H1127: READ <= 8'Hf2;
      32'H1128: READ <= 8'Hd8;
      32'H1129: READ <= 8'Ha4;
      32'H1130: READ <= 8'H8e;
      32'H1131: READ <= 8'H87;
      32'H1132: READ <= 8'H91;
      32'H1133: READ <= 8'H9d;
      32'H1134: READ <= 8'H9c;
      32'H1135: READ <= 8'Ha0;
      32'H1136: READ <= 8'H98;
      32'H1137: READ <= 8'Ha6;
      32'H1138: READ <= 8'H81;
      32'H1139: READ <= 8'H88;
      32'H1140: READ <= 8'H97;
      32'H1141: READ <= 8'H76;
      32'H1142: READ <= 8'H65;
      32'H1143: READ <= 8'H82;
      32'H1144: READ <= 8'H9e;
      32'H1145: READ <= 8'Ha8;
      32'H1146: READ <= 8'Had;
      32'H1147: READ <= 8'Hc3;
      32'H1148: READ <= 8'Hcd;
      32'H1149: READ <= 8'Hd0;
      32'H1150: READ <= 8'Hd1;
      32'H1151: READ <= 8'Hcb;
      32'H1152: READ <= 8'Hc3;
      32'H1153: READ <= 8'Hba;
      32'H1154: READ <= 8'Hc2;
      32'H1155: READ <= 8'Hcc;
      32'H1156: READ <= 8'Hca;
      32'H1157: READ <= 8'Hac;
      32'H1158: READ <= 8'H96;
      32'H1159: READ <= 8'Ha5;
      32'H1160: READ <= 8'H9b;
      32'H1161: READ <= 8'H98;
      32'H1162: READ <= 8'H92;
      32'H1163: READ <= 8'H8e;
      32'H1164: READ <= 8'H8e;
      32'H1165: READ <= 8'H8e;
      32'H1166: READ <= 8'H8e;
      32'H1167: READ <= 8'H8f;
      32'H1168: READ <= 8'H8e;
      32'H1169: READ <= 8'H8f;
      32'H1170: READ <= 8'H8f;
      32'H1171: READ <= 8'H90;
      32'H1172: READ <= 8'H91;
      32'H1173: READ <= 8'H91;
      32'H1174: READ <= 8'H91;
      32'H1175: READ <= 8'H92;
      32'H1176: READ <= 8'H93;
      32'H1177: READ <= 8'H95;
      32'H1178: READ <= 8'H96;
      32'H1179: READ <= 8'H96;
      32'H1180: READ <= 8'H97;
      32'H1181: READ <= 8'H97;
      32'H1182: READ <= 8'H97;
      32'H1183: READ <= 8'H98;
      32'H1184: READ <= 8'H97;
      32'H1185: READ <= 8'H98;
      32'H1186: READ <= 8'H98;
      32'H1187: READ <= 8'H98;
      32'H1188: READ <= 8'H99;
      32'H1189: READ <= 8'H99;
      32'H1190: READ <= 8'H99;
      32'H1191: READ <= 8'H99;
      32'H1192: READ <= 8'H9a;
      32'H1193: READ <= 8'H9a;
      32'H1194: READ <= 8'H9a;
      32'H1195: READ <= 8'H99;
      32'H1196: READ <= 8'H99;
      32'H1197: READ <= 8'H9a;
      32'H1198: READ <= 8'H9a;
      32'H1199: READ <= 8'H9b;
      32'H1200: READ <= 8'H9f;
      32'H1201: READ <= 8'Ha2;
      32'H1202: READ <= 8'Ha4;
      32'H1203: READ <= 8'Ha7;
      32'H1204: READ <= 8'Hab;
      32'H1205: READ <= 8'Hae;
      32'H1206: READ <= 8'Hb1;
      32'H1207: READ <= 8'Hb3;
      32'H1208: READ <= 8'Hb7;
      32'H1209: READ <= 8'Hba;
      32'H1210: READ <= 8'Hbd;
      32'H1211: READ <= 8'Hc0;
      32'H1212: READ <= 8'Hc4;
      32'H1213: READ <= 8'Hc9;
      32'H1214: READ <= 8'Hcc;
      32'H1215: READ <= 8'Hce;
      32'H1216: READ <= 8'Hd2;
      32'H1217: READ <= 8'Hd6;
      32'H1218: READ <= 8'Hda;
      32'H1219: READ <= 8'Hdf;
      32'H1220: READ <= 8'He2;
      32'H1221: READ <= 8'He5;
      32'H1222: READ <= 8'He8;
      32'H1223: READ <= 8'Hea;
      32'H1224: READ <= 8'Hec;
      32'H1225: READ <= 8'Hee;
      32'H1226: READ <= 8'Hec;
      32'H1227: READ <= 8'Hd8;
      32'H1228: READ <= 8'Ha9;
      32'H1229: READ <= 8'H87;
      32'H1230: READ <= 8'H87;
      32'H1231: READ <= 8'H83;
      32'H1232: READ <= 8'H8c;
      32'H1233: READ <= 8'H9b;
      32'H1234: READ <= 8'H9a;
      32'H1235: READ <= 8'H9f;
      32'H1236: READ <= 8'Ha3;
      32'H1237: READ <= 8'H99;
      32'H1238: READ <= 8'Hab;
      32'H1239: READ <= 8'H9c;
      32'H1240: READ <= 8'H8b;
      32'H1241: READ <= 8'H5a;
      32'H1242: READ <= 8'H40;
      32'H1243: READ <= 8'H72;
      32'H1244: READ <= 8'Ha7;
      32'H1245: READ <= 8'Hb0;
      32'H1246: READ <= 8'Hc8;
      32'H1247: READ <= 8'Hd8;
      32'H1248: READ <= 8'Hd6;
      32'H1249: READ <= 8'Hc0;
      32'H1250: READ <= 8'Hb5;
      32'H1251: READ <= 8'Hb9;
      32'H1252: READ <= 8'Hc7;
      32'H1253: READ <= 8'Hd8;
      32'H1254: READ <= 8'Hd8;
      32'H1255: READ <= 8'Hda;
      32'H1256: READ <= 8'Hd3;
      32'H1257: READ <= 8'Hcf;
      32'H1258: READ <= 8'Hba;
      32'H1259: READ <= 8'H9c;
      32'H1260: READ <= 8'H9f;
      32'H1261: READ <= 8'H96;
      32'H1262: READ <= 8'H96;
      32'H1263: READ <= 8'H93;
      32'H1264: READ <= 8'H8d;
      32'H1265: READ <= 8'H8d;
      32'H1266: READ <= 8'H8d;
      32'H1267: READ <= 8'H8e;
      32'H1268: READ <= 8'H8d;
      32'H1269: READ <= 8'H8e;
      32'H1270: READ <= 8'H8f;
      32'H1271: READ <= 8'H8f;
      32'H1272: READ <= 8'H8f;
      32'H1273: READ <= 8'H90;
      32'H1274: READ <= 8'H91;
      32'H1275: READ <= 8'H91;
      32'H1276: READ <= 8'H92;
      32'H1277: READ <= 8'H93;
      32'H1278: READ <= 8'H96;
      32'H1279: READ <= 8'H96;
      32'H1280: READ <= 8'H96;
      32'H1281: READ <= 8'H96;
      32'H1282: READ <= 8'H97;
      32'H1283: READ <= 8'H97;
      32'H1284: READ <= 8'H97;
      32'H1285: READ <= 8'H97;
      32'H1286: READ <= 8'H97;
      32'H1287: READ <= 8'H97;
      32'H1288: READ <= 8'H97;
      32'H1289: READ <= 8'H97;
      32'H1290: READ <= 8'H98;
      32'H1291: READ <= 8'H98;
      32'H1292: READ <= 8'H99;
      32'H1293: READ <= 8'H99;
      32'H1294: READ <= 8'H99;
      32'H1295: READ <= 8'H98;
      32'H1296: READ <= 8'H99;
      32'H1297: READ <= 8'H99;
      32'H1298: READ <= 8'H99;
      32'H1299: READ <= 8'H9a;
      32'H1300: READ <= 8'H9e;
      32'H1301: READ <= 8'Ha0;
      32'H1302: READ <= 8'Ha2;
      32'H1303: READ <= 8'Ha5;
      32'H1304: READ <= 8'Haa;
      32'H1305: READ <= 8'Had;
      32'H1306: READ <= 8'Haf;
      32'H1307: READ <= 8'Hb2;
      32'H1308: READ <= 8'Hb5;
      32'H1309: READ <= 8'Hb8;
      32'H1310: READ <= 8'Hbb;
      32'H1311: READ <= 8'Hbe;
      32'H1312: READ <= 8'Hc1;
      32'H1313: READ <= 8'Hc6;
      32'H1314: READ <= 8'Hca;
      32'H1315: READ <= 8'Hcd;
      32'H1316: READ <= 8'Hcf;
      32'H1317: READ <= 8'Hd3;
      32'H1318: READ <= 8'Hd9;
      32'H1319: READ <= 8'Hdd;
      32'H1320: READ <= 8'He1;
      32'H1321: READ <= 8'He5;
      32'H1322: READ <= 8'He7;
      32'H1323: READ <= 8'He9;
      32'H1324: READ <= 8'Hec;
      32'H1325: READ <= 8'Hed;
      32'H1326: READ <= 8'Hd9;
      32'H1327: READ <= 8'Ha8;
      32'H1328: READ <= 8'H9e;
      32'H1329: READ <= 8'H8c;
      32'H1330: READ <= 8'H82;
      32'H1331: READ <= 8'H89;
      32'H1332: READ <= 8'H95;
      32'H1333: READ <= 8'H95;
      32'H1334: READ <= 8'H99;
      32'H1335: READ <= 8'H90;
      32'H1336: READ <= 8'H9c;
      32'H1337: READ <= 8'H93;
      32'H1338: READ <= 8'H92;
      32'H1339: READ <= 8'H73;
      32'H1340: READ <= 8'H5a;
      32'H1341: READ <= 8'H2d;
      32'H1342: READ <= 8'H20;
      32'H1343: READ <= 8'H67;
      32'H1344: READ <= 8'Ha4;
      32'H1345: READ <= 8'Hbd;
      32'H1346: READ <= 8'Hcf;
      32'H1347: READ <= 8'Hbd;
      32'H1348: READ <= 8'Hab;
      32'H1349: READ <= 8'Hb0;
      32'H1350: READ <= 8'Hc4;
      32'H1351: READ <= 8'Hd9;
      32'H1352: READ <= 8'Hd5;
      32'H1353: READ <= 8'Hdd;
      32'H1354: READ <= 8'Hdd;
      32'H1355: READ <= 8'Hd7;
      32'H1356: READ <= 8'Hce;
      32'H1357: READ <= 8'Hc1;
      32'H1358: READ <= 8'Hba;
      32'H1359: READ <= 8'Haf;
      32'H1360: READ <= 8'Ha5;
      32'H1361: READ <= 8'H97;
      32'H1362: READ <= 8'H8d;
      32'H1363: READ <= 8'H8e;
      32'H1364: READ <= 8'H95;
      32'H1365: READ <= 8'H93;
      32'H1366: READ <= 8'H8d;
      32'H1367: READ <= 8'H8c;
      32'H1368: READ <= 8'H8d;
      32'H1369: READ <= 8'H8c;
      32'H1370: READ <= 8'H8d;
      32'H1371: READ <= 8'H8e;
      32'H1372: READ <= 8'H8e;
      32'H1373: READ <= 8'H8f;
      32'H1374: READ <= 8'H90;
      32'H1375: READ <= 8'H91;
      32'H1376: READ <= 8'H91;
      32'H1377: READ <= 8'H93;
      32'H1378: READ <= 8'H94;
      32'H1379: READ <= 8'H94;
      32'H1380: READ <= 8'H95;
      32'H1381: READ <= 8'H96;
      32'H1382: READ <= 8'H96;
      32'H1383: READ <= 8'H96;
      32'H1384: READ <= 8'H95;
      32'H1385: READ <= 8'H96;
      32'H1386: READ <= 8'H96;
      32'H1387: READ <= 8'H96;
      32'H1388: READ <= 8'H96;
      32'H1389: READ <= 8'H97;
      32'H1390: READ <= 8'H97;
      32'H1391: READ <= 8'H98;
      32'H1392: READ <= 8'H97;
      32'H1393: READ <= 8'H97;
      32'H1394: READ <= 8'H97;
      32'H1395: READ <= 8'H97;
      32'H1396: READ <= 8'H98;
      32'H1397: READ <= 8'H98;
      32'H1398: READ <= 8'H99;
      32'H1399: READ <= 8'H99;
      32'H1400: READ <= 8'H9e;
      32'H1401: READ <= 8'H9e;
      32'H1402: READ <= 8'Ha1;
      32'H1403: READ <= 8'Ha4;
      32'H1404: READ <= 8'Ha7;
      32'H1405: READ <= 8'Hab;
      32'H1406: READ <= 8'Hae;
      32'H1407: READ <= 8'Hb0;
      32'H1408: READ <= 8'Hb2;
      32'H1409: READ <= 8'Hb6;
      32'H1410: READ <= 8'Hb9;
      32'H1411: READ <= 8'Hbc;
      32'H1412: READ <= 8'Hc0;
      32'H1413: READ <= 8'Hc4;
      32'H1414: READ <= 8'Hc8;
      32'H1415: READ <= 8'Hcb;
      32'H1416: READ <= 8'Hcd;
      32'H1417: READ <= 8'Hd0;
      32'H1418: READ <= 8'Hd5;
      32'H1419: READ <= 8'Hda;
      32'H1420: READ <= 8'He0;
      32'H1421: READ <= 8'He3;
      32'H1422: READ <= 8'He7;
      32'H1423: READ <= 8'He9;
      32'H1424: READ <= 8'Hec;
      32'H1425: READ <= 8'He8;
      32'H1426: READ <= 8'Hc0;
      32'H1427: READ <= 8'H99;
      32'H1428: READ <= 8'H95;
      32'H1429: READ <= 8'H82;
      32'H1430: READ <= 8'H92;
      32'H1431: READ <= 8'H93;
      32'H1432: READ <= 8'Ha0;
      32'H1433: READ <= 8'H97;
      32'H1434: READ <= 8'H94;
      32'H1435: READ <= 8'H94;
      32'H1436: READ <= 8'H8f;
      32'H1437: READ <= 8'H7f;
      32'H1438: READ <= 8'H70;
      32'H1439: READ <= 8'H2e;
      32'H1440: READ <= 8'H14;
      32'H1441: READ <= 8'H1a;
      32'H1442: READ <= 8'H41;
      32'H1443: READ <= 8'H8c;
      32'H1444: READ <= 8'H8f;
      32'H1445: READ <= 8'H97;
      32'H1446: READ <= 8'H97;
      32'H1447: READ <= 8'Ha2;
      32'H1448: READ <= 8'Hb8;
      32'H1449: READ <= 8'Hd0;
      32'H1450: READ <= 8'Hda;
      32'H1451: READ <= 8'He2;
      32'H1452: READ <= 8'Hd9;
      32'H1453: READ <= 8'Hc7;
      32'H1454: READ <= 8'Hbe;
      32'H1455: READ <= 8'Hc1;
      32'H1456: READ <= 8'Hca;
      32'H1457: READ <= 8'Hcc;
      32'H1458: READ <= 8'Hd1;
      32'H1459: READ <= 8'Hd4;
      32'H1460: READ <= 8'Hd0;
      32'H1461: READ <= 8'Hd0;
      32'H1462: READ <= 8'Had;
      32'H1463: READ <= 8'H9d;
      32'H1464: READ <= 8'H9b;
      32'H1465: READ <= 8'H93;
      32'H1466: READ <= 8'H95;
      32'H1467: READ <= 8'H8e;
      32'H1468: READ <= 8'H8a;
      32'H1469: READ <= 8'H8b;
      32'H1470: READ <= 8'H8b;
      32'H1471: READ <= 8'H8c;
      32'H1472: READ <= 8'H8d;
      32'H1473: READ <= 8'H8e;
      32'H1474: READ <= 8'H8f;
      32'H1475: READ <= 8'H8f;
      32'H1476: READ <= 8'H8f;
      32'H1477: READ <= 8'H91;
      32'H1478: READ <= 8'H92;
      32'H1479: READ <= 8'H92;
      32'H1480: READ <= 8'H94;
      32'H1481: READ <= 8'H94;
      32'H1482: READ <= 8'H94;
      32'H1483: READ <= 8'H94;
      32'H1484: READ <= 8'H95;
      32'H1485: READ <= 8'H96;
      32'H1486: READ <= 8'H95;
      32'H1487: READ <= 8'H95;
      32'H1488: READ <= 8'H96;
      32'H1489: READ <= 8'H96;
      32'H1490: READ <= 8'H96;
      32'H1491: READ <= 8'H96;
      32'H1492: READ <= 8'H96;
      32'H1493: READ <= 8'H97;
      32'H1494: READ <= 8'H97;
      32'H1495: READ <= 8'H96;
      32'H1496: READ <= 8'H97;
      32'H1497: READ <= 8'H97;
      32'H1498: READ <= 8'H97;
      32'H1499: READ <= 8'H97;
      32'H1500: READ <= 8'H9c;
      32'H1501: READ <= 8'H9d;
      32'H1502: READ <= 8'Ha0;
      32'H1503: READ <= 8'Ha3;
      32'H1504: READ <= 8'Ha5;
      32'H1505: READ <= 8'Ha9;
      32'H1506: READ <= 8'Hac;
      32'H1507: READ <= 8'Haf;
      32'H1508: READ <= 8'Hb1;
      32'H1509: READ <= 8'Hb4;
      32'H1510: READ <= 8'Hb8;
      32'H1511: READ <= 8'Hbb;
      32'H1512: READ <= 8'Hbe;
      32'H1513: READ <= 8'Hc2;
      32'H1514: READ <= 8'Hc5;
      32'H1515: READ <= 8'Hc9;
      32'H1516: READ <= 8'Hcb;
      32'H1517: READ <= 8'Hcf;
      32'H1518: READ <= 8'Hd3;
      32'H1519: READ <= 8'Hd8;
      32'H1520: READ <= 8'Hdd;
      32'H1521: READ <= 8'He1;
      32'H1522: READ <= 8'He5;
      32'H1523: READ <= 8'Hea;
      32'H1524: READ <= 8'He9;
      32'H1525: READ <= 8'Hd2;
      32'H1526: READ <= 8'Haf;
      32'H1527: READ <= 8'Hab;
      32'H1528: READ <= 8'H98;
      32'H1529: READ <= 8'H89;
      32'H1530: READ <= 8'H92;
      32'H1531: READ <= 8'H90;
      32'H1532: READ <= 8'H98;
      32'H1533: READ <= 8'H89;
      32'H1534: READ <= 8'H7d;
      32'H1535: READ <= 8'H72;
      32'H1536: READ <= 8'H8a;
      32'H1537: READ <= 8'H62;
      32'H1538: READ <= 8'H34;
      32'H1539: READ <= 8'H1;
      32'H1540: READ <= 8'H16;
      32'H1541: READ <= 8'H5f;
      32'H1542: READ <= 8'H91;
      32'H1543: READ <= 8'Ha8;
      32'H1544: READ <= 8'H8f;
      32'H1545: READ <= 8'H82;
      32'H1546: READ <= 8'H9f;
      32'H1547: READ <= 8'Hcb;
      32'H1548: READ <= 8'Hcd;
      32'H1549: READ <= 8'Hc8;
      32'H1550: READ <= 8'Hbe;
      32'H1551: READ <= 8'Haf;
      32'H1552: READ <= 8'Had;
      32'H1553: READ <= 8'Hb3;
      32'H1554: READ <= 8'Hcf;
      32'H1555: READ <= 8'Hd9;
      32'H1556: READ <= 8'Hdc;
      32'H1557: READ <= 8'Hdf;
      32'H1558: READ <= 8'He8;
      32'H1559: READ <= 8'He7;
      32'H1560: READ <= 8'He0;
      32'H1561: READ <= 8'Hdd;
      32'H1562: READ <= 8'Hd7;
      32'H1563: READ <= 8'H9e;
      32'H1564: READ <= 8'H9a;
      32'H1565: READ <= 8'H91;
      32'H1566: READ <= 8'H87;
      32'H1567: READ <= 8'H8a;
      32'H1568: READ <= 8'H92;
      32'H1569: READ <= 8'H89;
      32'H1570: READ <= 8'H8a;
      32'H1571: READ <= 8'H8b;
      32'H1572: READ <= 8'H8c;
      32'H1573: READ <= 8'H8c;
      32'H1574: READ <= 8'H8e;
      32'H1575: READ <= 8'H8e;
      32'H1576: READ <= 8'H8f;
      32'H1577: READ <= 8'H8f;
      32'H1578: READ <= 8'H91;
      32'H1579: READ <= 8'H91;
      32'H1580: READ <= 8'H92;
      32'H1581: READ <= 8'H93;
      32'H1582: READ <= 8'H93;
      32'H1583: READ <= 8'H93;
      32'H1584: READ <= 8'H94;
      32'H1585: READ <= 8'H94;
      32'H1586: READ <= 8'H94;
      32'H1587: READ <= 8'H94;
      32'H1588: READ <= 8'H94;
      32'H1589: READ <= 8'H94;
      32'H1590: READ <= 8'H94;
      32'H1591: READ <= 8'H95;
      32'H1592: READ <= 8'H96;
      32'H1593: READ <= 8'H96;
      32'H1594: READ <= 8'H96;
      32'H1595: READ <= 8'H96;
      32'H1596: READ <= 8'H96;
      32'H1597: READ <= 8'H96;
      32'H1598: READ <= 8'H96;
      32'H1599: READ <= 8'H96;
      32'H1600: READ <= 8'H9a;
      32'H1601: READ <= 8'H9c;
      32'H1602: READ <= 8'H9e;
      32'H1603: READ <= 8'Ha0;
      32'H1604: READ <= 8'Ha4;
      32'H1605: READ <= 8'Ha7;
      32'H1606: READ <= 8'Haa;
      32'H1607: READ <= 8'Had;
      32'H1608: READ <= 8'Hb0;
      32'H1609: READ <= 8'Hb2;
      32'H1610: READ <= 8'Hb7;
      32'H1611: READ <= 8'Hba;
      32'H1612: READ <= 8'Hbc;
      32'H1613: READ <= 8'Hbe;
      32'H1614: READ <= 8'Hc3;
      32'H1615: READ <= 8'Hc7;
      32'H1616: READ <= 8'Hc9;
      32'H1617: READ <= 8'Hcd;
      32'H1618: READ <= 8'Hd0;
      32'H1619: READ <= 8'Hd6;
      32'H1620: READ <= 8'Hdb;
      32'H1621: READ <= 8'He0;
      32'H1622: READ <= 8'He3;
      32'H1623: READ <= 8'He6;
      32'H1624: READ <= 8'He9;
      32'H1625: READ <= 8'Hc7;
      32'H1626: READ <= 8'Haf;
      32'H1627: READ <= 8'Hb1;
      32'H1628: READ <= 8'H91;
      32'H1629: READ <= 8'H8d;
      32'H1630: READ <= 8'H9d;
      32'H1631: READ <= 8'H97;
      32'H1632: READ <= 8'H96;
      32'H1633: READ <= 8'H6d;
      32'H1634: READ <= 8'H82;
      32'H1635: READ <= 8'H6f;
      32'H1636: READ <= 8'H70;
      32'H1637: READ <= 8'H41;
      32'H1638: READ <= 8'H0;
      32'H1639: READ <= 8'H38;
      32'H1640: READ <= 8'H8c;
      32'H1641: READ <= 8'H97;
      32'H1642: READ <= 8'Ha8;
      32'H1643: READ <= 8'H88;
      32'H1644: READ <= 8'H86;
      32'H1645: READ <= 8'Hb3;
      32'H1646: READ <= 8'Hbd;
      32'H1647: READ <= 8'Hc3;
      32'H1648: READ <= 8'Hb0;
      32'H1649: READ <= 8'Had;
      32'H1650: READ <= 8'Haa;
      32'H1651: READ <= 8'Hb7;
      32'H1652: READ <= 8'Hc8;
      32'H1653: READ <= 8'Hd2;
      32'H1654: READ <= 8'Hd8;
      32'H1655: READ <= 8'Hd8;
      32'H1656: READ <= 8'Hdc;
      32'H1657: READ <= 8'He1;
      32'H1658: READ <= 8'He8;
      32'H1659: READ <= 8'Heb;
      32'H1660: READ <= 8'He7;
      32'H1661: READ <= 8'Hd9;
      32'H1662: READ <= 8'Hd5;
      32'H1663: READ <= 8'Hc2;
      32'H1664: READ <= 8'H86;
      32'H1665: READ <= 8'H82;
      32'H1666: READ <= 8'H82;
      32'H1667: READ <= 8'H7d;
      32'H1668: READ <= 8'H88;
      32'H1669: READ <= 8'H96;
      32'H1670: READ <= 8'H8c;
      32'H1671: READ <= 8'H8a;
      32'H1672: READ <= 8'H8a;
      32'H1673: READ <= 8'H8b;
      32'H1674: READ <= 8'H8c;
      32'H1675: READ <= 8'H8d;
      32'H1676: READ <= 8'H8d;
      32'H1677: READ <= 8'H8f;
      32'H1678: READ <= 8'H8f;
      32'H1679: READ <= 8'H90;
      32'H1680: READ <= 8'H91;
      32'H1681: READ <= 8'H92;
      32'H1682: READ <= 8'H92;
      32'H1683: READ <= 8'H92;
      32'H1684: READ <= 8'H93;
      32'H1685: READ <= 8'H92;
      32'H1686: READ <= 8'H92;
      32'H1687: READ <= 8'H93;
      32'H1688: READ <= 8'H93;
      32'H1689: READ <= 8'H93;
      32'H1690: READ <= 8'H94;
      32'H1691: READ <= 8'H94;
      32'H1692: READ <= 8'H94;
      32'H1693: READ <= 8'H95;
      32'H1694: READ <= 8'H95;
      32'H1695: READ <= 8'H95;
      32'H1696: READ <= 8'H95;
      32'H1697: READ <= 8'H95;
      32'H1698: READ <= 8'H95;
      32'H1699: READ <= 8'H95;
      32'H1700: READ <= 8'H97;
      32'H1701: READ <= 8'H9a;
      32'H1702: READ <= 8'H9b;
      32'H1703: READ <= 8'H9e;
      32'H1704: READ <= 8'Ha1;
      32'H1705: READ <= 8'Ha5;
      32'H1706: READ <= 8'Ha8;
      32'H1707: READ <= 8'Hab;
      32'H1708: READ <= 8'Hae;
      32'H1709: READ <= 8'Hb1;
      32'H1710: READ <= 8'Hb4;
      32'H1711: READ <= 8'Hb8;
      32'H1712: READ <= 8'Hbb;
      32'H1713: READ <= 8'Hbc;
      32'H1714: READ <= 8'Hc1;
      32'H1715: READ <= 8'Hc5;
      32'H1716: READ <= 8'Hc7;
      32'H1717: READ <= 8'Hca;
      32'H1718: READ <= 8'Hcf;
      32'H1719: READ <= 8'Hd4;
      32'H1720: READ <= 8'Hd8;
      32'H1721: READ <= 8'Hdd;
      32'H1722: READ <= 8'He1;
      32'H1723: READ <= 8'He4;
      32'H1724: READ <= 8'He2;
      32'H1725: READ <= 8'Hb1;
      32'H1726: READ <= 8'Hab;
      32'H1727: READ <= 8'Ha0;
      32'H1728: READ <= 8'H88;
      32'H1729: READ <= 8'H8f;
      32'H1730: READ <= 8'H9a;
      32'H1731: READ <= 8'H84;
      32'H1732: READ <= 8'H77;
      32'H1733: READ <= 8'H7a;
      32'H1734: READ <= 8'H71;
      32'H1735: READ <= 8'H73;
      32'H1736: READ <= 8'H57;
      32'H1737: READ <= 8'H26;
      32'H1738: READ <= 8'H2a;
      32'H1739: READ <= 8'H7e;
      32'H1740: READ <= 8'H79;
      32'H1741: READ <= 8'H8e;
      32'H1742: READ <= 8'Ha2;
      32'H1743: READ <= 8'H7f;
      32'H1744: READ <= 8'H63;
      32'H1745: READ <= 8'H80;
      32'H1746: READ <= 8'H9d;
      32'H1747: READ <= 8'H7c;
      32'H1748: READ <= 8'H85;
      32'H1749: READ <= 8'H91;
      32'H1750: READ <= 8'Ha3;
      32'H1751: READ <= 8'Ha4;
      32'H1752: READ <= 8'Haa;
      32'H1753: READ <= 8'Hb0;
      32'H1754: READ <= 8'Hb6;
      32'H1755: READ <= 8'Hb4;
      32'H1756: READ <= 8'Hb8;
      32'H1757: READ <= 8'Hc0;
      32'H1758: READ <= 8'Hc6;
      32'H1759: READ <= 8'Hce;
      32'H1760: READ <= 8'Hc7;
      32'H1761: READ <= 8'Hbc;
      32'H1762: READ <= 8'Hbe;
      32'H1763: READ <= 8'Hcd;
      32'H1764: READ <= 8'Hc5;
      32'H1765: READ <= 8'H9c;
      32'H1766: READ <= 8'H7f;
      32'H1767: READ <= 8'H8c;
      32'H1768: READ <= 8'H75;
      32'H1769: READ <= 8'H83;
      32'H1770: READ <= 8'H93;
      32'H1771: READ <= 8'H8e;
      32'H1772: READ <= 8'H88;
      32'H1773: READ <= 8'H89;
      32'H1774: READ <= 8'H8b;
      32'H1775: READ <= 8'H8b;
      32'H1776: READ <= 8'H8c;
      32'H1777: READ <= 8'H8d;
      32'H1778: READ <= 8'H8e;
      32'H1779: READ <= 8'H8f;
      32'H1780: READ <= 8'H8f;
      32'H1781: READ <= 8'H90;
      32'H1782: READ <= 8'H92;
      32'H1783: READ <= 8'H92;
      32'H1784: READ <= 8'H92;
      32'H1785: READ <= 8'H91;
      32'H1786: READ <= 8'H91;
      32'H1787: READ <= 8'H92;
      32'H1788: READ <= 8'H93;
      32'H1789: READ <= 8'H93;
      32'H1790: READ <= 8'H93;
      32'H1791: READ <= 8'H94;
      32'H1792: READ <= 8'H93;
      32'H1793: READ <= 8'H94;
      32'H1794: READ <= 8'H94;
      32'H1795: READ <= 8'H94;
      32'H1796: READ <= 8'H95;
      32'H1797: READ <= 8'H94;
      32'H1798: READ <= 8'H94;
      32'H1799: READ <= 8'H95;
      32'H1800: READ <= 8'H95;
      32'H1801: READ <= 8'H97;
      32'H1802: READ <= 8'H99;
      32'H1803: READ <= 8'H9b;
      32'H1804: READ <= 8'H9f;
      32'H1805: READ <= 8'Ha3;
      32'H1806: READ <= 8'Ha6;
      32'H1807: READ <= 8'Ha9;
      32'H1808: READ <= 8'Hac;
      32'H1809: READ <= 8'Haf;
      32'H1810: READ <= 8'Hb3;
      32'H1811: READ <= 8'Hb6;
      32'H1812: READ <= 8'Hb9;
      32'H1813: READ <= 8'Hbb;
      32'H1814: READ <= 8'Hbf;
      32'H1815: READ <= 8'Hc3;
      32'H1816: READ <= 8'Hc5;
      32'H1817: READ <= 8'Hc8;
      32'H1818: READ <= 8'Hcc;
      32'H1819: READ <= 8'Hd0;
      32'H1820: READ <= 8'Hd5;
      32'H1821: READ <= 8'Hdb;
      32'H1822: READ <= 8'Hde;
      32'H1823: READ <= 8'He1;
      32'H1824: READ <= 8'Hca;
      32'H1825: READ <= 8'Ha9;
      32'H1826: READ <= 8'Ha3;
      32'H1827: READ <= 8'H9e;
      32'H1828: READ <= 8'H7c;
      32'H1829: READ <= 8'H7e;
      32'H1830: READ <= 8'H7b;
      32'H1831: READ <= 8'H87;
      32'H1832: READ <= 8'H6c;
      32'H1833: READ <= 8'H82;
      32'H1834: READ <= 8'H82;
      32'H1835: READ <= 8'H74;
      32'H1836: READ <= 8'H5b;
      32'H1837: READ <= 8'Ha;
      32'H1838: READ <= 8'H4e;
      32'H1839: READ <= 8'H50;
      32'H1840: READ <= 8'H43;
      32'H1841: READ <= 8'H4d;
      32'H1842: READ <= 8'H71;
      32'H1843: READ <= 8'H63;
      32'H1844: READ <= 8'H6d;
      32'H1845: READ <= 8'H3d;
      32'H1846: READ <= 8'H5e;
      32'H1847: READ <= 8'H76;
      32'H1848: READ <= 8'H72;
      32'H1849: READ <= 8'H70;
      32'H1850: READ <= 8'H6c;
      32'H1851: READ <= 8'H6e;
      32'H1852: READ <= 8'H69;
      32'H1853: READ <= 8'H62;
      32'H1854: READ <= 8'H61;
      32'H1855: READ <= 8'H64;
      32'H1856: READ <= 8'H69;
      32'H1857: READ <= 8'H6e;
      32'H1858: READ <= 8'H7a;
      32'H1859: READ <= 8'H90;
      32'H1860: READ <= 8'H90;
      32'H1861: READ <= 8'H95;
      32'H1862: READ <= 8'H95;
      32'H1863: READ <= 8'H93;
      32'H1864: READ <= 8'H99;
      32'H1865: READ <= 8'H9c;
      32'H1866: READ <= 8'H9c;
      32'H1867: READ <= 8'H94;
      32'H1868: READ <= 8'H76;
      32'H1869: READ <= 8'H72;
      32'H1870: READ <= 8'H7b;
      32'H1871: READ <= 8'H8e;
      32'H1872: READ <= 8'H93;
      32'H1873: READ <= 8'H8a;
      32'H1874: READ <= 8'H8a;
      32'H1875: READ <= 8'H8a;
      32'H1876: READ <= 8'H8c;
      32'H1877: READ <= 8'H8c;
      32'H1878: READ <= 8'H8d;
      32'H1879: READ <= 8'H8e;
      32'H1880: READ <= 8'H8e;
      32'H1881: READ <= 8'H8f;
      32'H1882: READ <= 8'H8f;
      32'H1883: READ <= 8'H90;
      32'H1884: READ <= 8'H91;
      32'H1885: READ <= 8'H90;
      32'H1886: READ <= 8'H90;
      32'H1887: READ <= 8'H90;
      32'H1888: READ <= 8'H92;
      32'H1889: READ <= 8'H93;
      32'H1890: READ <= 8'H92;
      32'H1891: READ <= 8'H93;
      32'H1892: READ <= 8'H93;
      32'H1893: READ <= 8'H93;
      32'H1894: READ <= 8'H93;
      32'H1895: READ <= 8'H94;
      32'H1896: READ <= 8'H94;
      32'H1897: READ <= 8'H93;
      32'H1898: READ <= 8'H94;
      32'H1899: READ <= 8'H94;
      32'H1900: READ <= 8'H93;
      32'H1901: READ <= 8'H94;
      32'H1902: READ <= 8'H97;
      32'H1903: READ <= 8'H99;
      32'H1904: READ <= 8'H9c;
      32'H1905: READ <= 8'Ha0;
      32'H1906: READ <= 8'Ha4;
      32'H1907: READ <= 8'Ha7;
      32'H1908: READ <= 8'Haa;
      32'H1909: READ <= 8'Hae;
      32'H1910: READ <= 8'Hb1;
      32'H1911: READ <= 8'Hb3;
      32'H1912: READ <= 8'Hb7;
      32'H1913: READ <= 8'Hbb;
      32'H1914: READ <= 8'Hbe;
      32'H1915: READ <= 8'Hc1;
      32'H1916: READ <= 8'Hc4;
      32'H1917: READ <= 8'Hc6;
      32'H1918: READ <= 8'Hca;
      32'H1919: READ <= 8'Hcd;
      32'H1920: READ <= 8'Hd2;
      32'H1921: READ <= 8'Hd7;
      32'H1922: READ <= 8'Hdd;
      32'H1923: READ <= 8'Hdd;
      32'H1924: READ <= 8'Hb4;
      32'H1925: READ <= 8'Ha7;
      32'H1926: READ <= 8'H9f;
      32'H1927: READ <= 8'H93;
      32'H1928: READ <= 8'H6c;
      32'H1929: READ <= 8'H7f;
      32'H1930: READ <= 8'H77;
      32'H1931: READ <= 8'H70;
      32'H1932: READ <= 8'H7d;
      32'H1933: READ <= 8'H7f;
      32'H1934: READ <= 8'H6d;
      32'H1935: READ <= 8'H76;
      32'H1936: READ <= 8'H40;
      32'H1937: READ <= 8'H17;
      32'H1938: READ <= 8'H4c;
      32'H1939: READ <= 8'H48;
      32'H1940: READ <= 8'H2f;
      32'H1941: READ <= 8'H31;
      32'H1942: READ <= 8'H3c;
      32'H1943: READ <= 8'H20;
      32'H1944: READ <= 8'H2c;
      32'H1945: READ <= 8'H44;
      32'H1946: READ <= 8'H4a;
      32'H1947: READ <= 8'H5e;
      32'H1948: READ <= 8'H63;
      32'H1949: READ <= 8'H5f;
      32'H1950: READ <= 8'H59;
      32'H1951: READ <= 8'H54;
      32'H1952: READ <= 8'H51;
      32'H1953: READ <= 8'H50;
      32'H1954: READ <= 8'H58;
      32'H1955: READ <= 8'H61;
      32'H1956: READ <= 8'H6f;
      32'H1957: READ <= 8'H81;
      32'H1958: READ <= 8'H8f;
      32'H1959: READ <= 8'H9b;
      32'H1960: READ <= 8'H98;
      32'H1961: READ <= 8'H96;
      32'H1962: READ <= 8'H96;
      32'H1963: READ <= 8'H9e;
      32'H1964: READ <= 8'H9d;
      32'H1965: READ <= 8'H8b;
      32'H1966: READ <= 8'H74;
      32'H1967: READ <= 8'H71;
      32'H1968: READ <= 8'H76;
      32'H1969: READ <= 8'H7f;
      32'H1970: READ <= 8'H80;
      32'H1971: READ <= 8'H7b;
      32'H1972: READ <= 8'H8a;
      32'H1973: READ <= 8'H97;
      32'H1974: READ <= 8'H8e;
      32'H1975: READ <= 8'H89;
      32'H1976: READ <= 8'H8a;
      32'H1977: READ <= 8'H8b;
      32'H1978: READ <= 8'H8c;
      32'H1979: READ <= 8'H8c;
      32'H1980: READ <= 8'H8d;
      32'H1981: READ <= 8'H8e;
      32'H1982: READ <= 8'H8f;
      32'H1983: READ <= 8'H8f;
      32'H1984: READ <= 8'H8f;
      32'H1985: READ <= 8'H8f;
      32'H1986: READ <= 8'H8f;
      32'H1987: READ <= 8'H90;
      32'H1988: READ <= 8'H91;
      32'H1989: READ <= 8'H91;
      32'H1990: READ <= 8'H92;
      32'H1991: READ <= 8'H92;
      32'H1992: READ <= 8'H92;
      32'H1993: READ <= 8'H92;
      32'H1994: READ <= 8'H93;
      32'H1995: READ <= 8'H93;
      32'H1996: READ <= 8'H93;
      32'H1997: READ <= 8'H93;
      32'H1998: READ <= 8'H93;
      32'H1999: READ <= 8'H93;
      32'H2000: READ <= 8'H91;
      32'H2001: READ <= 8'H93;
      32'H2002: READ <= 8'H95;
      32'H2003: READ <= 8'H97;
      32'H2004: READ <= 8'H9a;
      32'H2005: READ <= 8'H9d;
      32'H2006: READ <= 8'Ha1;
      32'H2007: READ <= 8'Ha5;
      32'H2008: READ <= 8'Haa;
      32'H2009: READ <= 8'Hac;
      32'H2010: READ <= 8'Haf;
      32'H2011: READ <= 8'Hb1;
      32'H2012: READ <= 8'Hb5;
      32'H2013: READ <= 8'Hba;
      32'H2014: READ <= 8'Hbc;
      32'H2015: READ <= 8'Hbf;
      32'H2016: READ <= 8'Hc2;
      32'H2017: READ <= 8'Hc4;
      32'H2018: READ <= 8'Hc8;
      32'H2019: READ <= 8'Hcb;
      32'H2020: READ <= 8'Hd0;
      32'H2021: READ <= 8'Hd5;
      32'H2022: READ <= 8'Hda;
      32'H2023: READ <= 8'Hcc;
      32'H2024: READ <= 8'Hb3;
      32'H2025: READ <= 8'Ha9;
      32'H2026: READ <= 8'H94;
      32'H2027: READ <= 8'H87;
      32'H2028: READ <= 8'H5d;
      32'H2029: READ <= 8'H7e;
      32'H2030: READ <= 8'H6e;
      32'H2031: READ <= 8'H70;
      32'H2032: READ <= 8'H72;
      32'H2033: READ <= 8'H71;
      32'H2034: READ <= 8'H84;
      32'H2035: READ <= 8'H7a;
      32'H2036: READ <= 8'H42;
      32'H2037: READ <= 8'H14;
      32'H2038: READ <= 8'H42;
      32'H2039: READ <= 8'H2c;
      32'H2040: READ <= 8'H23;
      32'H2041: READ <= 8'H31;
      32'H2042: READ <= 8'H25;
      32'H2043: READ <= 8'H19;
      32'H2044: READ <= 8'H24;
      32'H2045: READ <= 8'H21;
      32'H2046: READ <= 8'H1c;
      32'H2047: READ <= 8'H38;
      32'H2048: READ <= 8'H43;
      32'H2049: READ <= 8'H32;
      32'H2050: READ <= 8'H2b;
      32'H2051: READ <= 8'H31;
      32'H2052: READ <= 8'H41;
      32'H2053: READ <= 8'H3a;
      32'H2054: READ <= 8'H2f;
      32'H2055: READ <= 8'H36;
      32'H2056: READ <= 8'H3a;
      32'H2057: READ <= 8'H3f;
      32'H2058: READ <= 8'H48;
      32'H2059: READ <= 8'H48;
      32'H2060: READ <= 8'H54;
      32'H2061: READ <= 8'H4a;
      32'H2062: READ <= 8'H40;
      32'H2063: READ <= 8'H49;
      32'H2064: READ <= 8'H53;
      32'H2065: READ <= 8'H56;
      32'H2066: READ <= 8'H44;
      32'H2067: READ <= 8'H41;
      32'H2068: READ <= 8'H47;
      32'H2069: READ <= 8'H52;
      32'H2070: READ <= 8'H64;
      32'H2071: READ <= 8'H74;
      32'H2072: READ <= 8'H79;
      32'H2073: READ <= 8'H84;
      32'H2074: READ <= 8'H93;
      32'H2075: READ <= 8'H8e;
      32'H2076: READ <= 8'H89;
      32'H2077: READ <= 8'H89;
      32'H2078: READ <= 8'H8a;
      32'H2079: READ <= 8'H8b;
      32'H2080: READ <= 8'H8c;
      32'H2081: READ <= 8'H8d;
      32'H2082: READ <= 8'H8d;
      32'H2083: READ <= 8'H8e;
      32'H2084: READ <= 8'H8d;
      32'H2085: READ <= 8'H8d;
      32'H2086: READ <= 8'H8d;
      32'H2087: READ <= 8'H8e;
      32'H2088: READ <= 8'H8f;
      32'H2089: READ <= 8'H90;
      32'H2090: READ <= 8'H90;
      32'H2091: READ <= 8'H91;
      32'H2092: READ <= 8'H92;
      32'H2093: READ <= 8'H92;
      32'H2094: READ <= 8'H92;
      32'H2095: READ <= 8'H92;
      32'H2096: READ <= 8'H91;
      32'H2097: READ <= 8'H92;
      32'H2098: READ <= 8'H91;
      32'H2099: READ <= 8'H91;
      32'H2100: READ <= 8'H90;
      32'H2101: READ <= 8'H91;
      32'H2102: READ <= 8'H93;
      32'H2103: READ <= 8'H95;
      32'H2104: READ <= 8'H97;
      32'H2105: READ <= 8'H9a;
      32'H2106: READ <= 8'H9e;
      32'H2107: READ <= 8'Ha2;
      32'H2108: READ <= 8'Ha7;
      32'H2109: READ <= 8'Hab;
      32'H2110: READ <= 8'Had;
      32'H2111: READ <= 8'Hb0;
      32'H2112: READ <= 8'Hb4;
      32'H2113: READ <= 8'Hb7;
      32'H2114: READ <= 8'Hbb;
      32'H2115: READ <= 8'Hbd;
      32'H2116: READ <= 8'Hbf;
      32'H2117: READ <= 8'Hc2;
      32'H2118: READ <= 8'Hc5;
      32'H2119: READ <= 8'Hc8;
      32'H2120: READ <= 8'Hcd;
      32'H2121: READ <= 8'Hd2;
      32'H2122: READ <= 8'Hc8;
      32'H2123: READ <= 8'Had;
      32'H2124: READ <= 8'Haa;
      32'H2125: READ <= 8'H8f;
      32'H2126: READ <= 8'H7a;
      32'H2127: READ <= 8'H71;
      32'H2128: READ <= 8'H56;
      32'H2129: READ <= 8'H7a;
      32'H2130: READ <= 8'H75;
      32'H2131: READ <= 8'H71;
      32'H2132: READ <= 8'H65;
      32'H2133: READ <= 8'H70;
      32'H2134: READ <= 8'H7d;
      32'H2135: READ <= 8'H7c;
      32'H2136: READ <= 8'H42;
      32'H2137: READ <= 8'He;
      32'H2138: READ <= 8'H2b;
      32'H2139: READ <= 8'H2b;
      32'H2140: READ <= 8'H22;
      32'H2141: READ <= 8'H29;
      32'H2142: READ <= 8'H23;
      32'H2143: READ <= 8'H21;
      32'H2144: READ <= 8'H23;
      32'H2145: READ <= 8'H29;
      32'H2146: READ <= 8'H2e;
      32'H2147: READ <= 8'H18;
      32'H2148: READ <= 8'H20;
      32'H2149: READ <= 8'H38;
      32'H2150: READ <= 8'H43;
      32'H2151: READ <= 8'H69;
      32'H2152: READ <= 8'H77;
      32'H2153: READ <= 8'H6f;
      32'H2154: READ <= 8'H5a;
      32'H2155: READ <= 8'H30;
      32'H2156: READ <= 8'H3d;
      32'H2157: READ <= 8'H56;
      32'H2158: READ <= 8'H6a;
      32'H2159: READ <= 8'H73;
      32'H2160: READ <= 8'H72;
      32'H2161: READ <= 8'H59;
      32'H2162: READ <= 8'H2d;
      32'H2163: READ <= 8'H21;
      32'H2164: READ <= 8'H26;
      32'H2165: READ <= 8'H33;
      32'H2166: READ <= 8'H36;
      32'H2167: READ <= 8'H2a;
      32'H2168: READ <= 8'H18;
      32'H2169: READ <= 8'H26;
      32'H2170: READ <= 8'H3e;
      32'H2171: READ <= 8'H54;
      32'H2172: READ <= 8'H79;
      32'H2173: READ <= 8'H7b;
      32'H2174: READ <= 8'H75;
      32'H2175: READ <= 8'H7f;
      32'H2176: READ <= 8'H8c;
      32'H2177: READ <= 8'H8b;
      32'H2178: READ <= 8'H88;
      32'H2179: READ <= 8'H89;
      32'H2180: READ <= 8'H8a;
      32'H2181: READ <= 8'H8b;
      32'H2182: READ <= 8'H8c;
      32'H2183: READ <= 8'H8c;
      32'H2184: READ <= 8'H8c;
      32'H2185: READ <= 8'H8c;
      32'H2186: READ <= 8'H8d;
      32'H2187: READ <= 8'H8c;
      32'H2188: READ <= 8'H8e;
      32'H2189: READ <= 8'H8f;
      32'H2190: READ <= 8'H8e;
      32'H2191: READ <= 8'H90;
      32'H2192: READ <= 8'H90;
      32'H2193: READ <= 8'H90;
      32'H2194: READ <= 8'H90;
      32'H2195: READ <= 8'H91;
      32'H2196: READ <= 8'H90;
      32'H2197: READ <= 8'H91;
      32'H2198: READ <= 8'H90;
      32'H2199: READ <= 8'H8f;
      32'H2200: READ <= 8'H8e;
      32'H2201: READ <= 8'H90;
      32'H2202: READ <= 8'H91;
      32'H2203: READ <= 8'H92;
      32'H2204: READ <= 8'H95;
      32'H2205: READ <= 8'H97;
      32'H2206: READ <= 8'H9b;
      32'H2207: READ <= 8'Ha0;
      32'H2208: READ <= 8'Ha3;
      32'H2209: READ <= 8'Ha8;
      32'H2210: READ <= 8'Hac;
      32'H2211: READ <= 8'Hae;
      32'H2212: READ <= 8'Hb1;
      32'H2213: READ <= 8'Hb4;
      32'H2214: READ <= 8'Hb8;
      32'H2215: READ <= 8'Hbb;
      32'H2216: READ <= 8'Hbd;
      32'H2217: READ <= 8'Hbf;
      32'H2218: READ <= 8'Hc1;
      32'H2219: READ <= 8'Hc6;
      32'H2220: READ <= 8'Hcd;
      32'H2221: READ <= 8'Hcc;
      32'H2222: READ <= 8'Hb1;
      32'H2223: READ <= 8'Ha3;
      32'H2224: READ <= 8'H9f;
      32'H2225: READ <= 8'H8d;
      32'H2226: READ <= 8'H6d;
      32'H2227: READ <= 8'H5e;
      32'H2228: READ <= 8'H42;
      32'H2229: READ <= 8'H68;
      32'H2230: READ <= 8'H79;
      32'H2231: READ <= 8'H7b;
      32'H2232: READ <= 8'H5a;
      32'H2233: READ <= 8'H3c;
      32'H2234: READ <= 8'H3e;
      32'H2235: READ <= 8'H35;
      32'H2236: READ <= 8'H29;
      32'H2237: READ <= 8'H23;
      32'H2238: READ <= 8'H1e;
      32'H2239: READ <= 8'H1b;
      32'H2240: READ <= 8'H13;
      32'H2241: READ <= 8'H1d;
      32'H2242: READ <= 8'H29;
      32'H2243: READ <= 8'H20;
      32'H2244: READ <= 8'H3c;
      32'H2245: READ <= 8'H40;
      32'H2246: READ <= 8'H3f;
      32'H2247: READ <= 8'H37;
      32'H2248: READ <= 8'H5a;
      32'H2249: READ <= 8'H72;
      32'H2250: READ <= 8'H72;
      32'H2251: READ <= 8'H6f;
      32'H2252: READ <= 8'H7a;
      32'H2253: READ <= 8'H70;
      32'H2254: READ <= 8'H63;
      32'H2255: READ <= 8'H14;
      32'H2256: READ <= 8'H14;
      32'H2257: READ <= 8'H20;
      32'H2258: READ <= 8'H34;
      32'H2259: READ <= 8'H51;
      32'H2260: READ <= 8'H62;
      32'H2261: READ <= 8'H73;
      32'H2262: READ <= 8'H46;
      32'H2263: READ <= 8'H38;
      32'H2264: READ <= 8'H6d;
      32'H2265: READ <= 8'H3a;
      32'H2266: READ <= 8'H3c;
      32'H2267: READ <= 8'H3b;
      32'H2268: READ <= 8'H2d;
      32'H2269: READ <= 8'H1f;
      32'H2270: READ <= 8'H1f;
      32'H2271: READ <= 8'H37;
      32'H2272: READ <= 8'H53;
      32'H2273: READ <= 8'H74;
      32'H2274: READ <= 8'H82;
      32'H2275: READ <= 8'H77;
      32'H2276: READ <= 8'H78;
      32'H2277: READ <= 8'H83;
      32'H2278: READ <= 8'H8a;
      32'H2279: READ <= 8'H88;
      32'H2280: READ <= 8'H89;
      32'H2281: READ <= 8'H89;
      32'H2282: READ <= 8'H8a;
      32'H2283: READ <= 8'H8a;
      32'H2284: READ <= 8'H8a;
      32'H2285: READ <= 8'H8b;
      32'H2286: READ <= 8'H8c;
      32'H2287: READ <= 8'H8b;
      32'H2288: READ <= 8'H8c;
      32'H2289: READ <= 8'H8d;
      32'H2290: READ <= 8'H8e;
      32'H2291: READ <= 8'H8e;
      32'H2292: READ <= 8'H8f;
      32'H2293: READ <= 8'H8e;
      32'H2294: READ <= 8'H8f;
      32'H2295: READ <= 8'H8f;
      32'H2296: READ <= 8'H8f;
      32'H2297: READ <= 8'H8f;
      32'H2298: READ <= 8'H8e;
      32'H2299: READ <= 8'H8e;
      32'H2300: READ <= 8'H8e;
      32'H2301: READ <= 8'H8e;
      32'H2302: READ <= 8'H8e;
      32'H2303: READ <= 8'H8f;
      32'H2304: READ <= 8'H91;
      32'H2305: READ <= 8'H94;
      32'H2306: READ <= 8'H98;
      32'H2307: READ <= 8'H9d;
      32'H2308: READ <= 8'Ha1;
      32'H2309: READ <= 8'Ha5;
      32'H2310: READ <= 8'Ha9;
      32'H2311: READ <= 8'Hac;
      32'H2312: READ <= 8'Hae;
      32'H2313: READ <= 8'Hb2;
      32'H2314: READ <= 8'Hb6;
      32'H2315: READ <= 8'Hb9;
      32'H2316: READ <= 8'Hba;
      32'H2317: READ <= 8'Hbc;
      32'H2318: READ <= 8'Hbf;
      32'H2319: READ <= 8'Hc3;
      32'H2320: READ <= 8'Hcb;
      32'H2321: READ <= 8'Hc7;
      32'H2322: READ <= 8'Haa;
      32'H2323: READ <= 8'H99;
      32'H2324: READ <= 8'H9a;
      32'H2325: READ <= 8'H99;
      32'H2326: READ <= 8'H8d;
      32'H2327: READ <= 8'H73;
      32'H2328: READ <= 8'H53;
      32'H2329: READ <= 8'H3f;
      32'H2330: READ <= 8'H5e;
      32'H2331: READ <= 8'H74;
      32'H2332: READ <= 8'H55;
      32'H2333: READ <= 8'H14;
      32'H2334: READ <= 8'He;
      32'H2335: READ <= 8'H12;
      32'H2336: READ <= 8'H14;
      32'H2337: READ <= 8'H3c;
      32'H2338: READ <= 8'H5b;
      32'H2339: READ <= 8'H50;
      32'H2340: READ <= 8'H45;
      32'H2341: READ <= 8'H34;
      32'H2342: READ <= 8'H1e;
      32'H2343: READ <= 8'H3;
      32'H2344: READ <= 8'H47;
      32'H2345: READ <= 8'H44;
      32'H2346: READ <= 8'H32;
      32'H2347: READ <= 8'H4c;
      32'H2348: READ <= 8'H69;
      32'H2349: READ <= 8'H6a;
      32'H2350: READ <= 8'H7a;
      32'H2351: READ <= 8'H78;
      32'H2352: READ <= 8'H6b;
      32'H2353: READ <= 8'H72;
      32'H2354: READ <= 8'H30;
      32'H2355: READ <= 8'H10;
      32'H2356: READ <= 8'H10;
      32'H2357: READ <= 8'H6;
      32'H2358: READ <= 8'H2;
      32'H2359: READ <= 8'Hd;
      32'H2360: READ <= 8'H16;
      32'H2361: READ <= 8'H41;
      32'H2362: READ <= 8'H50;
      32'H2363: READ <= 8'H44;
      32'H2364: READ <= 8'H82;
      32'H2365: READ <= 8'H52;
      32'H2366: READ <= 8'H66;
      32'H2367: READ <= 8'H65;
      32'H2368: READ <= 8'H68;
      32'H2369: READ <= 8'H4d;
      32'H2370: READ <= 8'H38;
      32'H2371: READ <= 8'H17;
      32'H2372: READ <= 8'H21;
      32'H2373: READ <= 8'H3f;
      32'H2374: READ <= 8'H6e;
      32'H2375: READ <= 8'H86;
      32'H2376: READ <= 8'H7a;
      32'H2377: READ <= 8'H74;
      32'H2378: READ <= 8'H7e;
      32'H2379: READ <= 8'H8a;
      32'H2380: READ <= 8'H87;
      32'H2381: READ <= 8'H89;
      32'H2382: READ <= 8'H89;
      32'H2383: READ <= 8'H89;
      32'H2384: READ <= 8'H8a;
      32'H2385: READ <= 8'H8a;
      32'H2386: READ <= 8'H8a;
      32'H2387: READ <= 8'H8a;
      32'H2388: READ <= 8'H8a;
      32'H2389: READ <= 8'H8c;
      32'H2390: READ <= 8'H8c;
      32'H2391: READ <= 8'H8c;
      32'H2392: READ <= 8'H8d;
      32'H2393: READ <= 8'H8d;
      32'H2394: READ <= 8'H8e;
      32'H2395: READ <= 8'H8e;
      32'H2396: READ <= 8'H8d;
      32'H2397: READ <= 8'H8d;
      32'H2398: READ <= 8'H8d;
      32'H2399: READ <= 8'H8c;
      32'H2400: READ <= 8'H8b;
      32'H2401: READ <= 8'H8b;
      32'H2402: READ <= 8'H8b;
      32'H2403: READ <= 8'H8c;
      32'H2404: READ <= 8'H8e;
      32'H2405: READ <= 8'H92;
      32'H2406: READ <= 8'H95;
      32'H2407: READ <= 8'H9a;
      32'H2408: READ <= 8'H9f;
      32'H2409: READ <= 8'Ha2;
      32'H2410: READ <= 8'Ha6;
      32'H2411: READ <= 8'Ha9;
      32'H2412: READ <= 8'Had;
      32'H2413: READ <= 8'Hb0;
      32'H2414: READ <= 8'Hb3;
      32'H2415: READ <= 8'Hb7;
      32'H2416: READ <= 8'Hb8;
      32'H2417: READ <= 8'Hba;
      32'H2418: READ <= 8'Hbc;
      32'H2419: READ <= 8'Hc2;
      32'H2420: READ <= 8'Hc5;
      32'H2421: READ <= 8'Hb3;
      32'H2422: READ <= 8'H9e;
      32'H2423: READ <= 8'H98;
      32'H2424: READ <= 8'H8e;
      32'H2425: READ <= 8'H8d;
      32'H2426: READ <= 8'H93;
      32'H2427: READ <= 8'H92;
      32'H2428: READ <= 8'H85;
      32'H2429: READ <= 8'H52;
      32'H2430: READ <= 8'H40;
      32'H2431: READ <= 8'H5f;
      32'H2432: READ <= 8'H54;
      32'H2433: READ <= 8'H5a;
      32'H2434: READ <= 8'H71;
      32'H2435: READ <= 8'H3e;
      32'H2436: READ <= 8'Ha;
      32'H2437: READ <= 8'H24;
      32'H2438: READ <= 8'H5f;
      32'H2439: READ <= 8'H62;
      32'H2440: READ <= 8'H59;
      32'H2441: READ <= 8'H80;
      32'H2442: READ <= 8'H5e;
      32'H2443: READ <= 8'H54;
      32'H2444: READ <= 8'H61;
      32'H2445: READ <= 8'H62;
      32'H2446: READ <= 8'H5d;
      32'H2447: READ <= 8'H4a;
      32'H2448: READ <= 8'H50;
      32'H2449: READ <= 8'H76;
      32'H2450: READ <= 8'H73;
      32'H2451: READ <= 8'H72;
      32'H2452: READ <= 8'H6c;
      32'H2453: READ <= 8'H60;
      32'H2454: READ <= 8'H3b;
      32'H2455: READ <= 8'H14;
      32'H2456: READ <= 8'H6;
      32'H2457: READ <= 8'H15;
      32'H2458: READ <= 8'H2b;
      32'H2459: READ <= 8'H14;
      32'H2460: READ <= 8'H4;
      32'H2461: READ <= 8'H2c;
      32'H2462: READ <= 8'H65;
      32'H2463: READ <= 8'H82;
      32'H2464: READ <= 8'H75;
      32'H2465: READ <= 8'H83;
      32'H2466: READ <= 8'Hb0;
      32'H2467: READ <= 8'Ha1;
      32'H2468: READ <= 8'Hac;
      32'H2469: READ <= 8'H9c;
      32'H2470: READ <= 8'H5f;
      32'H2471: READ <= 8'H4d;
      32'H2472: READ <= 8'H25;
      32'H2473: READ <= 8'H2a;
      32'H2474: READ <= 8'H36;
      32'H2475: READ <= 8'H56;
      32'H2476: READ <= 8'H72;
      32'H2477: READ <= 8'H84;
      32'H2478: READ <= 8'H78;
      32'H2479: READ <= 8'H78;
      32'H2480: READ <= 8'H89;
      32'H2481: READ <= 8'H87;
      32'H2482: READ <= 8'H88;
      32'H2483: READ <= 8'H88;
      32'H2484: READ <= 8'H89;
      32'H2485: READ <= 8'H8a;
      32'H2486: READ <= 8'H8a;
      32'H2487: READ <= 8'H8a;
      32'H2488: READ <= 8'H8a;
      32'H2489: READ <= 8'H8b;
      32'H2490: READ <= 8'H8b;
      32'H2491: READ <= 8'H8b;
      32'H2492: READ <= 8'H8c;
      32'H2493: READ <= 8'H8c;
      32'H2494: READ <= 8'H8c;
      32'H2495: READ <= 8'H8c;
      32'H2496: READ <= 8'H8b;
      32'H2497: READ <= 8'H8c;
      32'H2498: READ <= 8'H8b;
      32'H2499: READ <= 8'H8b;
      32'H2500: READ <= 8'H89;
      32'H2501: READ <= 8'H89;
      32'H2502: READ <= 8'H8a;
      32'H2503: READ <= 8'H8a;
      32'H2504: READ <= 8'H8c;
      32'H2505: READ <= 8'H8f;
      32'H2506: READ <= 8'H93;
      32'H2507: READ <= 8'H98;
      32'H2508: READ <= 8'H9d;
      32'H2509: READ <= 8'H9f;
      32'H2510: READ <= 8'Ha3;
      32'H2511: READ <= 8'Ha6;
      32'H2512: READ <= 8'Haa;
      32'H2513: READ <= 8'Had;
      32'H2514: READ <= 8'Hb1;
      32'H2515: READ <= 8'Hb3;
      32'H2516: READ <= 8'Hb6;
      32'H2517: READ <= 8'Hb8;
      32'H2518: READ <= 8'Hb9;
      32'H2519: READ <= 8'Hc1;
      32'H2520: READ <= 8'Hc9;
      32'H2521: READ <= 8'Ha7;
      32'H2522: READ <= 8'H88;
      32'H2523: READ <= 8'H88;
      32'H2524: READ <= 8'H8d;
      32'H2525: READ <= 8'H88;
      32'H2526: READ <= 8'H8b;
      32'H2527: READ <= 8'H90;
      32'H2528: READ <= 8'H96;
      32'H2529: READ <= 8'H94;
      32'H2530: READ <= 8'H8e;
      32'H2531: READ <= 8'H94;
      32'H2532: READ <= 8'H8c;
      32'H2533: READ <= 8'H97;
      32'H2534: READ <= 8'H97;
      32'H2535: READ <= 8'H81;
      32'H2536: READ <= 8'H58;
      32'H2537: READ <= 8'H20;
      32'H2538: READ <= 8'H42;
      32'H2539: READ <= 8'H5d;
      32'H2540: READ <= 8'H79;
      32'H2541: READ <= 8'H7d;
      32'H2542: READ <= 8'H8c;
      32'H2543: READ <= 8'H87;
      32'H2544: READ <= 8'H70;
      32'H2545: READ <= 8'H75;
      32'H2546: READ <= 8'H5b;
      32'H2547: READ <= 8'H5c;
      32'H2548: READ <= 8'H5a;
      32'H2549: READ <= 8'H41;
      32'H2550: READ <= 8'H78;
      32'H2551: READ <= 8'H75;
      32'H2552: READ <= 8'H4d;
      32'H2553: READ <= 8'H29;
      32'H2554: READ <= 8'H48;
      32'H2555: READ <= 8'Hc;
      32'H2556: READ <= 8'H9;
      32'H2557: READ <= 8'H26;
      32'H2558: READ <= 8'H4a;
      32'H2559: READ <= 8'H6f;
      32'H2560: READ <= 8'H6;
      32'H2561: READ <= 8'Ha;
      32'H2562: READ <= 8'H5b;
      32'H2563: READ <= 8'Ha3;
      32'H2564: READ <= 8'H9c;
      32'H2565: READ <= 8'Haa;
      32'H2566: READ <= 8'Hb7;
      32'H2567: READ <= 8'Hc1;
      32'H2568: READ <= 8'Hc0;
      32'H2569: READ <= 8'Hbf;
      32'H2570: READ <= 8'Ha3;
      32'H2571: READ <= 8'H6f;
      32'H2572: READ <= 8'H73;
      32'H2573: READ <= 8'H36;
      32'H2574: READ <= 8'H30;
      32'H2575: READ <= 8'H51;
      32'H2576: READ <= 8'H3a;
      32'H2577: READ <= 8'H41;
      32'H2578: READ <= 8'H74;
      32'H2579: READ <= 8'H8d;
      32'H2580: READ <= 8'H7b;
      32'H2581: READ <= 8'H88;
      32'H2582: READ <= 8'H88;
      32'H2583: READ <= 8'H88;
      32'H2584: READ <= 8'H88;
      32'H2585: READ <= 8'H88;
      32'H2586: READ <= 8'H89;
      32'H2587: READ <= 8'H89;
      32'H2588: READ <= 8'H89;
      32'H2589: READ <= 8'H89;
      32'H2590: READ <= 8'H89;
      32'H2591: READ <= 8'H8a;
      32'H2592: READ <= 8'H8a;
      32'H2593: READ <= 8'H8a;
      32'H2594: READ <= 8'H8a;
      32'H2595: READ <= 8'H8a;
      32'H2596: READ <= 8'H8b;
      32'H2597: READ <= 8'H8b;
      32'H2598: READ <= 8'H8a;
      32'H2599: READ <= 8'H8a;
      32'H2600: READ <= 8'H87;
      32'H2601: READ <= 8'H87;
      32'H2602: READ <= 8'H89;
      32'H2603: READ <= 8'H89;
      32'H2604: READ <= 8'H8a;
      32'H2605: READ <= 8'H8c;
      32'H2606: READ <= 8'H91;
      32'H2607: READ <= 8'H95;
      32'H2608: READ <= 8'H99;
      32'H2609: READ <= 8'H9d;
      32'H2610: READ <= 8'H9f;
      32'H2611: READ <= 8'Ha3;
      32'H2612: READ <= 8'Ha7;
      32'H2613: READ <= 8'Hab;
      32'H2614: READ <= 8'Haf;
      32'H2615: READ <= 8'Hb2;
      32'H2616: READ <= 8'Hb4;
      32'H2617: READ <= 8'Hb5;
      32'H2618: READ <= 8'Hb7;
      32'H2619: READ <= 8'Hc1;
      32'H2620: READ <= 8'Hc3;
      32'H2621: READ <= 8'H99;
      32'H2622: READ <= 8'H80;
      32'H2623: READ <= 8'H85;
      32'H2624: READ <= 8'H7f;
      32'H2625: READ <= 8'H85;
      32'H2626: READ <= 8'H86;
      32'H2627: READ <= 8'H86;
      32'H2628: READ <= 8'H8e;
      32'H2629: READ <= 8'H8f;
      32'H2630: READ <= 8'H90;
      32'H2631: READ <= 8'H8a;
      32'H2632: READ <= 8'H95;
      32'H2633: READ <= 8'H98;
      32'H2634: READ <= 8'H88;
      32'H2635: READ <= 8'H73;
      32'H2636: READ <= 8'H79;
      32'H2637: READ <= 8'H4d;
      32'H2638: READ <= 8'H5a;
      32'H2639: READ <= 8'H6b;
      32'H2640: READ <= 8'H81;
      32'H2641: READ <= 8'H7c;
      32'H2642: READ <= 8'H71;
      32'H2643: READ <= 8'H6f;
      32'H2644: READ <= 8'H6d;
      32'H2645: READ <= 8'H7d;
      32'H2646: READ <= 8'H79;
      32'H2647: READ <= 8'H66;
      32'H2648: READ <= 8'H55;
      32'H2649: READ <= 8'H3c;
      32'H2650: READ <= 8'H4e;
      32'H2651: READ <= 8'H47;
      32'H2652: READ <= 8'H10;
      32'H2653: READ <= 8'H32;
      32'H2654: READ <= 8'H43;
      32'H2655: READ <= 8'Hd;
      32'H2656: READ <= 8'H8;
      32'H2657: READ <= 8'H34;
      32'H2658: READ <= 8'H46;
      32'H2659: READ <= 8'H8f;
      32'H2660: READ <= 8'H35;
      32'H2661: READ <= 8'H0;
      32'H2662: READ <= 8'H49;
      32'H2663: READ <= 8'Hab;
      32'H2664: READ <= 8'Hb8;
      32'H2665: READ <= 8'Hbb;
      32'H2666: READ <= 8'Hba;
      32'H2667: READ <= 8'Hc1;
      32'H2668: READ <= 8'Hb7;
      32'H2669: READ <= 8'Hbd;
      32'H2670: READ <= 8'Hc5;
      32'H2671: READ <= 8'H93;
      32'H2672: READ <= 8'H87;
      32'H2673: READ <= 8'H80;
      32'H2674: READ <= 8'H6c;
      32'H2675: READ <= 8'H49;
      32'H2676: READ <= 8'H43;
      32'H2677: READ <= 8'H2b;
      32'H2678: READ <= 8'H28;
      32'H2679: READ <= 8'H4b;
      32'H2680: READ <= 8'H80;
      32'H2681: READ <= 8'H92;
      32'H2682: READ <= 8'H89;
      32'H2683: READ <= 8'H87;
      32'H2684: READ <= 8'H87;
      32'H2685: READ <= 8'H88;
      32'H2686: READ <= 8'H88;
      32'H2687: READ <= 8'H88;
      32'H2688: READ <= 8'H88;
      32'H2689: READ <= 8'H88;
      32'H2690: READ <= 8'H88;
      32'H2691: READ <= 8'H88;
      32'H2692: READ <= 8'H89;
      32'H2693: READ <= 8'H88;
      32'H2694: READ <= 8'H89;
      32'H2695: READ <= 8'H88;
      32'H2696: READ <= 8'H89;
      32'H2697: READ <= 8'H8a;
      32'H2698: READ <= 8'H8a;
      32'H2699: READ <= 8'H89;
      32'H2700: READ <= 8'H85;
      32'H2701: READ <= 8'H86;
      32'H2702: READ <= 8'H87;
      32'H2703: READ <= 8'H88;
      32'H2704: READ <= 8'H88;
      32'H2705: READ <= 8'H8b;
      32'H2706: READ <= 8'H8d;
      32'H2707: READ <= 8'H91;
      32'H2708: READ <= 8'H95;
      32'H2709: READ <= 8'H9a;
      32'H2710: READ <= 8'H9d;
      32'H2711: READ <= 8'Ha0;
      32'H2712: READ <= 8'Ha5;
      32'H2713: READ <= 8'Ha8;
      32'H2714: READ <= 8'Hac;
      32'H2715: READ <= 8'Hb0;
      32'H2716: READ <= 8'Hb1;
      32'H2717: READ <= 8'Hb3;
      32'H2718: READ <= 8'Hb6;
      32'H2719: READ <= 8'Hc0;
      32'H2720: READ <= 8'Hc2;
      32'H2721: READ <= 8'H92;
      32'H2722: READ <= 8'H89;
      32'H2723: READ <= 8'H89;
      32'H2724: READ <= 8'H76;
      32'H2725: READ <= 8'H7b;
      32'H2726: READ <= 8'H78;
      32'H2727: READ <= 8'H7b;
      32'H2728: READ <= 8'H8d;
      32'H2729: READ <= 8'H8a;
      32'H2730: READ <= 8'H8d;
      32'H2731: READ <= 8'H80;
      32'H2732: READ <= 8'H76;
      32'H2733: READ <= 8'H7a;
      32'H2734: READ <= 8'H80;
      32'H2735: READ <= 8'H72;
      32'H2736: READ <= 8'H75;
      32'H2737: READ <= 8'H34;
      32'H2738: READ <= 8'H49;
      32'H2739: READ <= 8'H6b;
      32'H2740: READ <= 8'H52;
      32'H2741: READ <= 8'H55;
      32'H2742: READ <= 8'H68;
      32'H2743: READ <= 8'H70;
      32'H2744: READ <= 8'H6f;
      32'H2745: READ <= 8'H61;
      32'H2746: READ <= 8'H74;
      32'H2747: READ <= 8'H6f;
      32'H2748: READ <= 8'H4e;
      32'H2749: READ <= 8'H4c;
      32'H2750: READ <= 8'H24;
      32'H2751: READ <= 8'H7;
      32'H2752: READ <= 8'H1a;
      32'H2753: READ <= 8'H43;
      32'H2754: READ <= 8'H49;
      32'H2755: READ <= 8'H9;
      32'H2756: READ <= 8'H6;
      32'H2757: READ <= 8'H18;
      32'H2758: READ <= 8'H62;
      32'H2759: READ <= 8'H94;
      32'H2760: READ <= 8'Haf;
      32'H2761: READ <= 8'H5;
      32'H2762: READ <= 8'H31;
      32'H2763: READ <= 8'Ha3;
      32'H2764: READ <= 8'H9d;
      32'H2765: READ <= 8'Hb2;
      32'H2766: READ <= 8'Hb6;
      32'H2767: READ <= 8'Hba;
      32'H2768: READ <= 8'Hbf;
      32'H2769: READ <= 8'Hc1;
      32'H2770: READ <= 8'Hbf;
      32'H2771: READ <= 8'Hb3;
      32'H2772: READ <= 8'H84;
      32'H2773: READ <= 8'H94;
      32'H2774: READ <= 8'H93;
      32'H2775: READ <= 8'H8d;
      32'H2776: READ <= 8'H74;
      32'H2777: READ <= 8'H84;
      32'H2778: READ <= 8'H51;
      32'H2779: READ <= 8'H38;
      32'H2780: READ <= 8'H32;
      32'H2781: READ <= 8'H5b;
      32'H2782: READ <= 8'H7d;
      32'H2783: READ <= 8'H87;
      32'H2784: READ <= 8'H86;
      32'H2785: READ <= 8'H87;
      32'H2786: READ <= 8'H87;
      32'H2787: READ <= 8'H87;
      32'H2788: READ <= 8'H88;
      32'H2789: READ <= 8'H87;
      32'H2790: READ <= 8'H87;
      32'H2791: READ <= 8'H88;
      32'H2792: READ <= 8'H88;
      32'H2793: READ <= 8'H87;
      32'H2794: READ <= 8'H88;
      32'H2795: READ <= 8'H88;
      32'H2796: READ <= 8'H88;
      32'H2797: READ <= 8'H88;
      32'H2798: READ <= 8'H89;
      32'H2799: READ <= 8'H89;
      32'H2800: READ <= 8'H83;
      32'H2801: READ <= 8'H84;
      32'H2802: READ <= 8'H85;
      32'H2803: READ <= 8'H87;
      32'H2804: READ <= 8'H87;
      32'H2805: READ <= 8'H89;
      32'H2806: READ <= 8'H8c;
      32'H2807: READ <= 8'H8f;
      32'H2808: READ <= 8'H93;
      32'H2809: READ <= 8'H97;
      32'H2810: READ <= 8'H9b;
      32'H2811: READ <= 8'H9e;
      32'H2812: READ <= 8'Ha3;
      32'H2813: READ <= 8'Ha5;
      32'H2814: READ <= 8'Ha9;
      32'H2815: READ <= 8'Hac;
      32'H2816: READ <= 8'Haf;
      32'H2817: READ <= 8'Hb0;
      32'H2818: READ <= 8'Hb3;
      32'H2819: READ <= 8'Hbe;
      32'H2820: READ <= 8'Hc5;
      32'H2821: READ <= 8'Ha0;
      32'H2822: READ <= 8'H91;
      32'H2823: READ <= 8'H78;
      32'H2824: READ <= 8'H7e;
      32'H2825: READ <= 8'H74;
      32'H2826: READ <= 8'H72;
      32'H2827: READ <= 8'H82;
      32'H2828: READ <= 8'H77;
      32'H2829: READ <= 8'H8b;
      32'H2830: READ <= 8'H7b;
      32'H2831: READ <= 8'H85;
      32'H2832: READ <= 8'H76;
      32'H2833: READ <= 8'H80;
      32'H2834: READ <= 8'H62;
      32'H2835: READ <= 8'H56;
      32'H2836: READ <= 8'H16;
      32'H2837: READ <= 8'H14;
      32'H2838: READ <= 8'H45;
      32'H2839: READ <= 8'H6b;
      32'H2840: READ <= 8'H65;
      32'H2841: READ <= 8'H68;
      32'H2842: READ <= 8'H65;
      32'H2843: READ <= 8'H61;
      32'H2844: READ <= 8'H5f;
      32'H2845: READ <= 8'H69;
      32'H2846: READ <= 8'H72;
      32'H2847: READ <= 8'H8a;
      32'H2848: READ <= 8'H5d;
      32'H2849: READ <= 8'H4e;
      32'H2850: READ <= 8'H22;
      32'H2851: READ <= 8'H1;
      32'H2852: READ <= 8'H22;
      32'H2853: READ <= 8'H53;
      32'H2854: READ <= 8'H49;
      32'H2855: READ <= 8'H9;
      32'H2856: READ <= 8'H6;
      32'H2857: READ <= 8'H1b;
      32'H2858: READ <= 8'H67;
      32'H2859: READ <= 8'H85;
      32'H2860: READ <= 8'Hb4;
      32'H2861: READ <= 8'H45;
      32'H2862: READ <= 8'H1b;
      32'H2863: READ <= 8'H9f;
      32'H2864: READ <= 8'Hb6;
      32'H2865: READ <= 8'Ha8;
      32'H2866: READ <= 8'Hb1;
      32'H2867: READ <= 8'Hb4;
      32'H2868: READ <= 8'Hb7;
      32'H2869: READ <= 8'Hbf;
      32'H2870: READ <= 8'Hc2;
      32'H2871: READ <= 8'Hb9;
      32'H2872: READ <= 8'H8b;
      32'H2873: READ <= 8'H65;
      32'H2874: READ <= 8'H8c;
      32'H2875: READ <= 8'Ha4;
      32'H2876: READ <= 8'Ha0;
      32'H2877: READ <= 8'Ha0;
      32'H2878: READ <= 8'H9a;
      32'H2879: READ <= 8'H54;
      32'H2880: READ <= 8'H49;
      32'H2881: READ <= 8'H47;
      32'H2882: READ <= 8'H40;
      32'H2883: READ <= 8'H58;
      32'H2884: READ <= 8'H85;
      32'H2885: READ <= 8'H87;
      32'H2886: READ <= 8'H86;
      32'H2887: READ <= 8'H86;
      32'H2888: READ <= 8'H86;
      32'H2889: READ <= 8'H86;
      32'H2890: READ <= 8'H86;
      32'H2891: READ <= 8'H87;
      32'H2892: READ <= 8'H87;
      32'H2893: READ <= 8'H86;
      32'H2894: READ <= 8'H88;
      32'H2895: READ <= 8'H87;
      32'H2896: READ <= 8'H87;
      32'H2897: READ <= 8'H88;
      32'H2898: READ <= 8'H88;
      32'H2899: READ <= 8'H89;
      32'H2900: READ <= 8'H83;
      32'H2901: READ <= 8'H83;
      32'H2902: READ <= 8'H84;
      32'H2903: READ <= 8'H84;
      32'H2904: READ <= 8'H85;
      32'H2905: READ <= 8'H87;
      32'H2906: READ <= 8'H89;
      32'H2907: READ <= 8'H8b;
      32'H2908: READ <= 8'H90;
      32'H2909: READ <= 8'H93;
      32'H2910: READ <= 8'H98;
      32'H2911: READ <= 8'H9b;
      32'H2912: READ <= 8'Ha0;
      32'H2913: READ <= 8'Ha3;
      32'H2914: READ <= 8'Ha6;
      32'H2915: READ <= 8'Ha8;
      32'H2916: READ <= 8'Hac;
      32'H2917: READ <= 8'Hae;
      32'H2918: READ <= 8'Hb2;
      32'H2919: READ <= 8'Hbb;
      32'H2920: READ <= 8'Hc1;
      32'H2921: READ <= 8'H9e;
      32'H2922: READ <= 8'H82;
      32'H2923: READ <= 8'H84;
      32'H2924: READ <= 8'H79;
      32'H2925: READ <= 8'H74;
      32'H2926: READ <= 8'H73;
      32'H2927: READ <= 8'H7d;
      32'H2928: READ <= 8'H7b;
      32'H2929: READ <= 8'H8c;
      32'H2930: READ <= 8'H84;
      32'H2931: READ <= 8'H7d;
      32'H2932: READ <= 8'H70;
      32'H2933: READ <= 8'H6a;
      32'H2934: READ <= 8'H55;
      32'H2935: READ <= 8'H13;
      32'H2936: READ <= 8'H8;
      32'H2937: READ <= 8'H1b;
      32'H2938: READ <= 8'H44;
      32'H2939: READ <= 8'H5a;
      32'H2940: READ <= 8'H4d;
      32'H2941: READ <= 8'H51;
      32'H2942: READ <= 8'H59;
      32'H2943: READ <= 8'H5e;
      32'H2944: READ <= 8'H82;
      32'H2945: READ <= 8'H69;
      32'H2946: READ <= 8'H5c;
      32'H2947: READ <= 8'H5f;
      32'H2948: READ <= 8'H65;
      32'H2949: READ <= 8'H50;
      32'H2950: READ <= 8'H2b;
      32'H2951: READ <= 8'H15;
      32'H2952: READ <= 8'H32;
      32'H2953: READ <= 8'H61;
      32'H2954: READ <= 8'H43;
      32'H2955: READ <= 8'Hc;
      32'H2956: READ <= 8'Ha;
      32'H2957: READ <= 8'H1b;
      32'H2958: READ <= 8'H63;
      32'H2959: READ <= 8'H8c;
      32'H2960: READ <= 8'Ha0;
      32'H2961: READ <= 8'H6e;
      32'H2962: READ <= 8'Hb;
      32'H2963: READ <= 8'H76;
      32'H2964: READ <= 8'Ha4;
      32'H2965: READ <= 8'Haa;
      32'H2966: READ <= 8'Hac;
      32'H2967: READ <= 8'Hac;
      32'H2968: READ <= 8'Hb7;
      32'H2969: READ <= 8'Hba;
      32'H2970: READ <= 8'Hc0;
      32'H2971: READ <= 8'Hb9;
      32'H2972: READ <= 8'H97;
      32'H2973: READ <= 8'H4e;
      32'H2974: READ <= 8'H4f;
      32'H2975: READ <= 8'Ha4;
      32'H2976: READ <= 8'Hb0;
      32'H2977: READ <= 8'Ha6;
      32'H2978: READ <= 8'Ha9;
      32'H2979: READ <= 8'H99;
      32'H2980: READ <= 8'H7f;
      32'H2981: READ <= 8'H92;
      32'H2982: READ <= 8'H64;
      32'H2983: READ <= 8'H4c;
      32'H2984: READ <= 8'H5a;
      32'H2985: READ <= 8'H85;
      32'H2986: READ <= 8'H87;
      32'H2987: READ <= 8'H86;
      32'H2988: READ <= 8'H86;
      32'H2989: READ <= 8'H86;
      32'H2990: READ <= 8'H86;
      32'H2991: READ <= 8'H86;
      32'H2992: READ <= 8'H86;
      32'H2993: READ <= 8'H86;
      32'H2994: READ <= 8'H87;
      32'H2995: READ <= 8'H87;
      32'H2996: READ <= 8'H87;
      32'H2997: READ <= 8'H88;
      32'H2998: READ <= 8'H88;
      32'H2999: READ <= 8'H88;
      32'H3000: READ <= 8'H82;
      32'H3001: READ <= 8'H82;
      32'H3002: READ <= 8'H82;
      32'H3003: READ <= 8'H83;
      32'H3004: READ <= 8'H84;
      32'H3005: READ <= 8'H85;
      32'H3006: READ <= 8'H87;
      32'H3007: READ <= 8'H89;
      32'H3008: READ <= 8'H8d;
      32'H3009: READ <= 8'H90;
      32'H3010: READ <= 8'H95;
      32'H3011: READ <= 8'H99;
      32'H3012: READ <= 8'H9c;
      32'H3013: READ <= 8'H9f;
      32'H3014: READ <= 8'Ha2;
      32'H3015: READ <= 8'Ha5;
      32'H3016: READ <= 8'Ha9;
      32'H3017: READ <= 8'Hab;
      32'H3018: READ <= 8'Hac;
      32'H3019: READ <= 8'Hbb;
      32'H3020: READ <= 8'Hc9;
      32'H3021: READ <= 8'H99;
      32'H3022: READ <= 8'H83;
      32'H3023: READ <= 8'H78;
      32'H3024: READ <= 8'H71;
      32'H3025: READ <= 8'H6b;
      32'H3026: READ <= 8'H72;
      32'H3027: READ <= 8'H74;
      32'H3028: READ <= 8'H74;
      32'H3029: READ <= 8'H81;
      32'H3030: READ <= 8'H7d;
      32'H3031: READ <= 8'H75;
      32'H3032: READ <= 8'H6f;
      32'H3033: READ <= 8'H63;
      32'H3034: READ <= 8'H3b;
      32'H3035: READ <= 8'H20;
      32'H3036: READ <= 8'H13;
      32'H3037: READ <= 8'H6;
      32'H3038: READ <= 8'H3c;
      32'H3039: READ <= 8'H4f;
      32'H3040: READ <= 8'H51;
      32'H3041: READ <= 8'H4c;
      32'H3042: READ <= 8'H6c;
      32'H3043: READ <= 8'H6d;
      32'H3044: READ <= 8'H72;
      32'H3045: READ <= 8'H7d;
      32'H3046: READ <= 8'H6e;
      32'H3047: READ <= 8'H7c;
      32'H3048: READ <= 8'H4a;
      32'H3049: READ <= 8'H41;
      32'H3050: READ <= 8'H19;
      32'H3051: READ <= 8'H2b;
      32'H3052: READ <= 8'H31;
      32'H3053: READ <= 8'H60;
      32'H3054: READ <= 8'H3c;
      32'H3055: READ <= 8'H8;
      32'H3056: READ <= 8'H6;
      32'H3057: READ <= 8'H1a;
      32'H3058: READ <= 8'H63;
      32'H3059: READ <= 8'H82;
      32'H3060: READ <= 8'H8d;
      32'H3061: READ <= 8'H7a;
      32'H3062: READ <= 8'H0;
      32'H3063: READ <= 8'H63;
      32'H3064: READ <= 8'Ha1;
      32'H3065: READ <= 8'H9d;
      32'H3066: READ <= 8'H9b;
      32'H3067: READ <= 8'Ha5;
      32'H3068: READ <= 8'Haa;
      32'H3069: READ <= 8'Had;
      32'H3070: READ <= 8'Hb7;
      32'H3071: READ <= 8'Hb5;
      32'H3072: READ <= 8'H98;
      32'H3073: READ <= 8'H4f;
      32'H3074: READ <= 8'H39;
      32'H3075: READ <= 8'H69;
      32'H3076: READ <= 8'Ha8;
      32'H3077: READ <= 8'Hb4;
      32'H3078: READ <= 8'Had;
      32'H3079: READ <= 8'Ha0;
      32'H3080: READ <= 8'H97;
      32'H3081: READ <= 8'H95;
      32'H3082: READ <= 8'H92;
      32'H3083: READ <= 8'H6f;
      32'H3084: READ <= 8'H5a;
      32'H3085: READ <= 8'H67;
      32'H3086: READ <= 8'H89;
      32'H3087: READ <= 8'H85;
      32'H3088: READ <= 8'H85;
      32'H3089: READ <= 8'H85;
      32'H3090: READ <= 8'H84;
      32'H3091: READ <= 8'H85;
      32'H3092: READ <= 8'H85;
      32'H3093: READ <= 8'H86;
      32'H3094: READ <= 8'H86;
      32'H3095: READ <= 8'H87;
      32'H3096: READ <= 8'H87;
      32'H3097: READ <= 8'H87;
      32'H3098: READ <= 8'H88;
      32'H3099: READ <= 8'H88;
      32'H3100: READ <= 8'H81;
      32'H3101: READ <= 8'H81;
      32'H3102: READ <= 8'H81;
      32'H3103: READ <= 8'H81;
      32'H3104: READ <= 8'H82;
      32'H3105: READ <= 8'H83;
      32'H3106: READ <= 8'H84;
      32'H3107: READ <= 8'H86;
      32'H3108: READ <= 8'H8a;
      32'H3109: READ <= 8'H8e;
      32'H3110: READ <= 8'H91;
      32'H3111: READ <= 8'H95;
      32'H3112: READ <= 8'H99;
      32'H3113: READ <= 8'H9c;
      32'H3114: READ <= 8'H9f;
      32'H3115: READ <= 8'Ha1;
      32'H3116: READ <= 8'Ha5;
      32'H3117: READ <= 8'Ha8;
      32'H3118: READ <= 8'Haa;
      32'H3119: READ <= 8'Hb1;
      32'H3120: READ <= 8'Hc5;
      32'H3121: READ <= 8'Ha0;
      32'H3122: READ <= 8'H80;
      32'H3123: READ <= 8'H71;
      32'H3124: READ <= 8'H6a;
      32'H3125: READ <= 8'H77;
      32'H3126: READ <= 8'H77;
      32'H3127: READ <= 8'H77;
      32'H3128: READ <= 8'H6d;
      32'H3129: READ <= 8'H6f;
      32'H3130: READ <= 8'H76;
      32'H3131: READ <= 8'H74;
      32'H3132: READ <= 8'H59;
      32'H3133: READ <= 8'H51;
      32'H3134: READ <= 8'H35;
      32'H3135: READ <= 8'H33;
      32'H3136: READ <= 8'H9;
      32'H3137: READ <= 8'H1;
      32'H3138: READ <= 8'H9;
      32'H3139: READ <= 8'H4b;
      32'H3140: READ <= 8'H45;
      32'H3141: READ <= 8'H56;
      32'H3142: READ <= 8'H50;
      32'H3143: READ <= 8'H60;
      32'H3144: READ <= 8'H67;
      32'H3145: READ <= 8'H58;
      32'H3146: READ <= 8'H64;
      32'H3147: READ <= 8'H5a;
      32'H3148: READ <= 8'H63;
      32'H3149: READ <= 8'H51;
      32'H3150: READ <= 8'H1b;
      32'H3151: READ <= 8'H36;
      32'H3152: READ <= 8'H34;
      32'H3153: READ <= 8'H66;
      32'H3154: READ <= 8'H2e;
      32'H3155: READ <= 8'H5;
      32'H3156: READ <= 8'H6;
      32'H3157: READ <= 8'H21;
      32'H3158: READ <= 8'H6c;
      32'H3159: READ <= 8'H82;
      32'H3160: READ <= 8'H90;
      32'H3161: READ <= 8'H7e;
      32'H3162: READ <= 8'H1;
      32'H3163: READ <= 8'H28;
      32'H3164: READ <= 8'H9a;
      32'H3165: READ <= 8'Ha7;
      32'H3166: READ <= 8'H9f;
      32'H3167: READ <= 8'H9d;
      32'H3168: READ <= 8'Hab;
      32'H3169: READ <= 8'Ha7;
      32'H3170: READ <= 8'Haa;
      32'H3171: READ <= 8'Ha8;
      32'H3172: READ <= 8'H8f;
      32'H3173: READ <= 8'H54;
      32'H3174: READ <= 8'H5e;
      32'H3175: READ <= 8'H4d;
      32'H3176: READ <= 8'H6b;
      32'H3177: READ <= 8'Ha0;
      32'H3178: READ <= 8'Ha6;
      32'H3179: READ <= 8'Ha7;
      32'H3180: READ <= 8'H8f;
      32'H3181: READ <= 8'Ha3;
      32'H3182: READ <= 8'Ha4;
      32'H3183: READ <= 8'H91;
      32'H3184: READ <= 8'H73;
      32'H3185: READ <= 8'H63;
      32'H3186: READ <= 8'H6f;
      32'H3187: READ <= 8'H86;
      32'H3188: READ <= 8'H86;
      32'H3189: READ <= 8'H84;
      32'H3190: READ <= 8'H84;
      32'H3191: READ <= 8'H85;
      32'H3192: READ <= 8'H85;
      32'H3193: READ <= 8'H85;
      32'H3194: READ <= 8'H86;
      32'H3195: READ <= 8'H86;
      32'H3196: READ <= 8'H88;
      32'H3197: READ <= 8'H87;
      32'H3198: READ <= 8'H88;
      32'H3199: READ <= 8'H88;
      32'H3200: READ <= 8'H7f;
      32'H3201: READ <= 8'H80;
      32'H3202: READ <= 8'H80;
      32'H3203: READ <= 8'H80;
      32'H3204: READ <= 8'H80;
      32'H3205: READ <= 8'H81;
      32'H3206: READ <= 8'H82;
      32'H3207: READ <= 8'H84;
      32'H3208: READ <= 8'H87;
      32'H3209: READ <= 8'H89;
      32'H3210: READ <= 8'H8d;
      32'H3211: READ <= 8'H92;
      32'H3212: READ <= 8'H95;
      32'H3213: READ <= 8'H98;
      32'H3214: READ <= 8'H9c;
      32'H3215: READ <= 8'H9e;
      32'H3216: READ <= 8'Ha2;
      32'H3217: READ <= 8'Ha4;
      32'H3218: READ <= 8'Ha6;
      32'H3219: READ <= 8'Hba;
      32'H3220: READ <= 8'Hcf;
      32'H3221: READ <= 8'Ha2;
      32'H3222: READ <= 8'H7d;
      32'H3223: READ <= 8'H6b;
      32'H3224: READ <= 8'H6e;
      32'H3225: READ <= 8'H6d;
      32'H3226: READ <= 8'H74;
      32'H3227: READ <= 8'H6b;
      32'H3228: READ <= 8'H76;
      32'H3229: READ <= 8'H7e;
      32'H3230: READ <= 8'H6a;
      32'H3231: READ <= 8'H66;
      32'H3232: READ <= 8'H69;
      32'H3233: READ <= 8'H54;
      32'H3234: READ <= 8'H29;
      32'H3235: READ <= 8'H2d;
      32'H3236: READ <= 8'H7;
      32'H3237: READ <= 8'H7;
      32'H3238: READ <= 8'H2;
      32'H3239: READ <= 8'H3f;
      32'H3240: READ <= 8'H3f;
      32'H3241: READ <= 8'H51;
      32'H3242: READ <= 8'H59;
      32'H3243: READ <= 8'H4e;
      32'H3244: READ <= 8'H6a;
      32'H3245: READ <= 8'H67;
      32'H3246: READ <= 8'H65;
      32'H3247: READ <= 8'H58;
      32'H3248: READ <= 8'H46;
      32'H3249: READ <= 8'H55;
      32'H3250: READ <= 8'H1a;
      32'H3251: READ <= 8'H40;
      32'H3252: READ <= 8'H41;
      32'H3253: READ <= 8'H67;
      32'H3254: READ <= 8'H1f;
      32'H3255: READ <= 8'H3;
      32'H3256: READ <= 8'H5;
      32'H3257: READ <= 8'H28;
      32'H3258: READ <= 8'H74;
      32'H3259: READ <= 8'H7a;
      32'H3260: READ <= 8'H95;
      32'H3261: READ <= 8'H93;
      32'H3262: READ <= 8'H2;
      32'H3263: READ <= 8'H3;
      32'H3264: READ <= 8'H76;
      32'H3265: READ <= 8'H9a;
      32'H3266: READ <= 8'Ha2;
      32'H3267: READ <= 8'Ha5;
      32'H3268: READ <= 8'Ha1;
      32'H3269: READ <= 8'H9f;
      32'H3270: READ <= 8'H99;
      32'H3271: READ <= 8'H9a;
      32'H3272: READ <= 8'H81;
      32'H3273: READ <= 8'H71;
      32'H3274: READ <= 8'H72;
      32'H3275: READ <= 8'H70;
      32'H3276: READ <= 8'H48;
      32'H3277: READ <= 8'H77;
      32'H3278: READ <= 8'H8c;
      32'H3279: READ <= 8'Hac;
      32'H3280: READ <= 8'H9d;
      32'H3281: READ <= 8'H95;
      32'H3282: READ <= 8'Ha8;
      32'H3283: READ <= 8'Hab;
      32'H3284: READ <= 8'H94;
      32'H3285: READ <= 8'H73;
      32'H3286: READ <= 8'H68;
      32'H3287: READ <= 8'H72;
      32'H3288: READ <= 8'H80;
      32'H3289: READ <= 8'H87;
      32'H3290: READ <= 8'H84;
      32'H3291: READ <= 8'H85;
      32'H3292: READ <= 8'H85;
      32'H3293: READ <= 8'H86;
      32'H3294: READ <= 8'H86;
      32'H3295: READ <= 8'H87;
      32'H3296: READ <= 8'H87;
      32'H3297: READ <= 8'H88;
      32'H3298: READ <= 8'H88;
      32'H3299: READ <= 8'H88;
      32'H3300: READ <= 8'H7e;
      32'H3301: READ <= 8'H7e;
      32'H3302: READ <= 8'H7e;
      32'H3303: READ <= 8'H7f;
      32'H3304: READ <= 8'H80;
      32'H3305: READ <= 8'H80;
      32'H3306: READ <= 8'H81;
      32'H3307: READ <= 8'H82;
      32'H3308: READ <= 8'H84;
      32'H3309: READ <= 8'H86;
      32'H3310: READ <= 8'H88;
      32'H3311: READ <= 8'H8d;
      32'H3312: READ <= 8'H90;
      32'H3313: READ <= 8'H93;
      32'H3314: READ <= 8'H97;
      32'H3315: READ <= 8'H9b;
      32'H3316: READ <= 8'H9e;
      32'H3317: READ <= 8'Ha3;
      32'H3318: READ <= 8'Hae;
      32'H3319: READ <= 8'Hc9;
      32'H3320: READ <= 8'Hcf;
      32'H3321: READ <= 8'H99;
      32'H3322: READ <= 8'H71;
      32'H3323: READ <= 8'H68;
      32'H3324: READ <= 8'H68;
      32'H3325: READ <= 8'H65;
      32'H3326: READ <= 8'H64;
      32'H3327: READ <= 8'H68;
      32'H3328: READ <= 8'H5d;
      32'H3329: READ <= 8'H57;
      32'H3330: READ <= 8'H5e;
      32'H3331: READ <= 8'H64;
      32'H3332: READ <= 8'H60;
      32'H3333: READ <= 8'H33;
      32'H3334: READ <= 8'H17;
      32'H3335: READ <= 8'H1d;
      32'H3336: READ <= 8'Hb;
      32'H3337: READ <= 8'Ha;
      32'H3338: READ <= 8'H4;
      32'H3339: READ <= 8'H8;
      32'H3340: READ <= 8'H49;
      32'H3341: READ <= 8'H4d;
      32'H3342: READ <= 8'H52;
      32'H3343: READ <= 8'H59;
      32'H3344: READ <= 8'H4d;
      32'H3345: READ <= 8'H6d;
      32'H3346: READ <= 8'H6e;
      32'H3347: READ <= 8'H57;
      32'H3348: READ <= 8'H63;
      32'H3349: READ <= 8'H4b;
      32'H3350: READ <= 8'H33;
      32'H3351: READ <= 8'H2c;
      32'H3352: READ <= 8'H4a;
      32'H3353: READ <= 8'H5f;
      32'H3354: READ <= 8'H1c;
      32'H3355: READ <= 8'H3;
      32'H3356: READ <= 8'H4;
      32'H3357: READ <= 8'H22;
      32'H3358: READ <= 8'H74;
      32'H3359: READ <= 8'H75;
      32'H3360: READ <= 8'H91;
      32'H3361: READ <= 8'H97;
      32'H3362: READ <= 8'H9;
      32'H3363: READ <= 8'H6;
      32'H3364: READ <= 8'H48;
      32'H3365: READ <= 8'Ha0;
      32'H3366: READ <= 8'H9b;
      32'H3367: READ <= 8'Ha0;
      32'H3368: READ <= 8'H9c;
      32'H3369: READ <= 8'H98;
      32'H3370: READ <= 8'H92;
      32'H3371: READ <= 8'H8d;
      32'H3372: READ <= 8'H90;
      32'H3373: READ <= 8'H94;
      32'H3374: READ <= 8'H89;
      32'H3375: READ <= 8'H7d;
      32'H3376: READ <= 8'H59;
      32'H3377: READ <= 8'H71;
      32'H3378: READ <= 8'H82;
      32'H3379: READ <= 8'H89;
      32'H3380: READ <= 8'H9c;
      32'H3381: READ <= 8'H90;
      32'H3382: READ <= 8'H9d;
      32'H3383: READ <= 8'Hb1;
      32'H3384: READ <= 8'Haf;
      32'H3385: READ <= 8'H8a;
      32'H3386: READ <= 8'H7c;
      32'H3387: READ <= 8'H6f;
      32'H3388: READ <= 8'H70;
      32'H3389: READ <= 8'H79;
      32'H3390: READ <= 8'H85;
      32'H3391: READ <= 8'H85;
      32'H3392: READ <= 8'H85;
      32'H3393: READ <= 8'H85;
      32'H3394: READ <= 8'H86;
      32'H3395: READ <= 8'H87;
      32'H3396: READ <= 8'H87;
      32'H3397: READ <= 8'H87;
      32'H3398: READ <= 8'H88;
      32'H3399: READ <= 8'H88;
      32'H3400: READ <= 8'H7c;
      32'H3401: READ <= 8'H7d;
      32'H3402: READ <= 8'H7d;
      32'H3403: READ <= 8'H7e;
      32'H3404: READ <= 8'H7e;
      32'H3405: READ <= 8'H7f;
      32'H3406: READ <= 8'H7f;
      32'H3407: READ <= 8'H81;
      32'H3408: READ <= 8'H81;
      32'H3409: READ <= 8'H84;
      32'H3410: READ <= 8'H85;
      32'H3411: READ <= 8'H86;
      32'H3412: READ <= 8'H8b;
      32'H3413: READ <= 8'H90;
      32'H3414: READ <= 8'H93;
      32'H3415: READ <= 8'H96;
      32'H3416: READ <= 8'H9a;
      32'H3417: READ <= 8'Ha2;
      32'H3418: READ <= 8'Hc2;
      32'H3419: READ <= 8'Hdd;
      32'H3420: READ <= 8'Hab;
      32'H3421: READ <= 8'H84;
      32'H3422: READ <= 8'H70;
      32'H3423: READ <= 8'H50;
      32'H3424: READ <= 8'H3b;
      32'H3425: READ <= 8'H35;
      32'H3426: READ <= 8'H33;
      32'H3427: READ <= 8'H51;
      32'H3428: READ <= 8'H51;
      32'H3429: READ <= 8'H5f;
      32'H3430: READ <= 8'H4b;
      32'H3431: READ <= 8'H45;
      32'H3432: READ <= 8'H47;
      32'H3433: READ <= 8'H3b;
      32'H3434: READ <= 8'H9;
      32'H3435: READ <= 8'H13;
      32'H3436: READ <= 8'H33;
      32'H3437: READ <= 8'H1f;
      32'H3438: READ <= 8'H10;
      32'H3439: READ <= 8'H7;
      32'H3440: READ <= 8'H15;
      32'H3441: READ <= 8'H44;
      32'H3442: READ <= 8'H3b;
      32'H3443: READ <= 8'H50;
      32'H3444: READ <= 8'H58;
      32'H3445: READ <= 8'H3e;
      32'H3446: READ <= 8'H54;
      32'H3447: READ <= 8'H50;
      32'H3448: READ <= 8'H71;
      32'H3449: READ <= 8'H2e;
      32'H3450: READ <= 8'H3e;
      32'H3451: READ <= 8'H2c;
      32'H3452: READ <= 8'H54;
      32'H3453: READ <= 8'H4f;
      32'H3454: READ <= 8'H17;
      32'H3455: READ <= 8'H4;
      32'H3456: READ <= 8'H3;
      32'H3457: READ <= 8'H1f;
      32'H3458: READ <= 8'H6e;
      32'H3459: READ <= 8'H7b;
      32'H3460: READ <= 8'H93;
      32'H3461: READ <= 8'H92;
      32'H3462: READ <= 8'He;
      32'H3463: READ <= 8'Hd;
      32'H3464: READ <= 8'H1c;
      32'H3465: READ <= 8'H94;
      32'H3466: READ <= 8'H98;
      32'H3467: READ <= 8'H91;
      32'H3468: READ <= 8'H93;
      32'H3469: READ <= 8'H8e;
      32'H3470: READ <= 8'H82;
      32'H3471: READ <= 8'H8a;
      32'H3472: READ <= 8'H91;
      32'H3473: READ <= 8'H9b;
      32'H3474: READ <= 8'H86;
      32'H3475: READ <= 8'H7d;
      32'H3476: READ <= 8'H5e;
      32'H3477: READ <= 8'H68;
      32'H3478: READ <= 8'H84;
      32'H3479: READ <= 8'H80;
      32'H3480: READ <= 8'H84;
      32'H3481: READ <= 8'H85;
      32'H3482: READ <= 8'H87;
      32'H3483: READ <= 8'H8d;
      32'H3484: READ <= 8'H94;
      32'H3485: READ <= 8'H85;
      32'H3486: READ <= 8'H92;
      32'H3487: READ <= 8'H87;
      32'H3488: READ <= 8'H84;
      32'H3489: READ <= 8'H7a;
      32'H3490: READ <= 8'H7c;
      32'H3491: READ <= 8'H85;
      32'H3492: READ <= 8'H85;
      32'H3493: READ <= 8'H86;
      32'H3494: READ <= 8'H87;
      32'H3495: READ <= 8'H87;
      32'H3496: READ <= 8'H87;
      32'H3497: READ <= 8'H88;
      32'H3498: READ <= 8'H88;
      32'H3499: READ <= 8'H88;
      32'H3500: READ <= 8'H7c;
      32'H3501: READ <= 8'H7c;
      32'H3502: READ <= 8'H7c;
      32'H3503: READ <= 8'H7c;
      32'H3504: READ <= 8'H7d;
      32'H3505: READ <= 8'H7d;
      32'H3506: READ <= 8'H7e;
      32'H3507: READ <= 8'H80;
      32'H3508: READ <= 8'H80;
      32'H3509: READ <= 8'H81;
      32'H3510: READ <= 8'H83;
      32'H3511: READ <= 8'H83;
      32'H3512: READ <= 8'H86;
      32'H3513: READ <= 8'H8a;
      32'H3514: READ <= 8'H8e;
      32'H3515: READ <= 8'H92;
      32'H3516: READ <= 8'H96;
      32'H3517: READ <= 8'Ha2;
      32'H3518: READ <= 8'Hc8;
      32'H3519: READ <= 8'Hb6;
      32'H3520: READ <= 8'H81;
      32'H3521: READ <= 8'H6c;
      32'H3522: READ <= 8'H6b;
      32'H3523: READ <= 8'H3d;
      32'H3524: READ <= 8'H20;
      32'H3525: READ <= 8'H16;
      32'H3526: READ <= 8'H13;
      32'H3527: READ <= 8'H12;
      32'H3528: READ <= 8'H17;
      32'H3529: READ <= 8'H1a;
      32'H3530: READ <= 8'H1f;
      32'H3531: READ <= 8'H46;
      32'H3532: READ <= 8'Hc;
      32'H3533: READ <= 8'H11;
      32'H3534: READ <= 8'H4;
      32'H3535: READ <= 8'H2b;
      32'H3536: READ <= 8'H37;
      32'H3537: READ <= 8'H3a;
      32'H3538: READ <= 8'H1e;
      32'H3539: READ <= 8'H7;
      32'H3540: READ <= 8'H7;
      32'H3541: READ <= 8'H2e;
      32'H3542: READ <= 8'H64;
      32'H3543: READ <= 8'H32;
      32'H3544: READ <= 8'H60;
      32'H3545: READ <= 8'H5a;
      32'H3546: READ <= 8'H4b;
      32'H3547: READ <= 8'H57;
      32'H3548: READ <= 8'H41;
      32'H3549: READ <= 8'H4e;
      32'H3550: READ <= 8'H3f;
      32'H3551: READ <= 8'H20;
      32'H3552: READ <= 8'H63;
      32'H3553: READ <= 8'H4e;
      32'H3554: READ <= 8'Hc;
      32'H3555: READ <= 8'H4;
      32'H3556: READ <= 8'Ha;
      32'H3557: READ <= 8'H23;
      32'H3558: READ <= 8'H6c;
      32'H3559: READ <= 8'H77;
      32'H3560: READ <= 8'H8d;
      32'H3561: READ <= 8'H97;
      32'H3562: READ <= 8'H19;
      32'H3563: READ <= 8'H1a;
      32'H3564: READ <= 8'Hf;
      32'H3565: READ <= 8'H77;
      32'H3566: READ <= 8'H8d;
      32'H3567: READ <= 8'H90;
      32'H3568: READ <= 8'H7f;
      32'H3569: READ <= 8'H76;
      32'H3570: READ <= 8'H7a;
      32'H3571: READ <= 8'H92;
      32'H3572: READ <= 8'H99;
      32'H3573: READ <= 8'H9e;
      32'H3574: READ <= 8'H8c;
      32'H3575: READ <= 8'H80;
      32'H3576: READ <= 8'H70;
      32'H3577: READ <= 8'H63;
      32'H3578: READ <= 8'H7e;
      32'H3579: READ <= 8'H7f;
      32'H3580: READ <= 8'H80;
      32'H3581: READ <= 8'H81;
      32'H3582: READ <= 8'H82;
      32'H3583: READ <= 8'H82;
      32'H3584: READ <= 8'H83;
      32'H3585: READ <= 8'H85;
      32'H3586: READ <= 8'H7a;
      32'H3587: READ <= 8'H79;
      32'H3588: READ <= 8'H8f;
      32'H3589: READ <= 8'H89;
      32'H3590: READ <= 8'H88;
      32'H3591: READ <= 8'H85;
      32'H3592: READ <= 8'H86;
      32'H3593: READ <= 8'H86;
      32'H3594: READ <= 8'H87;
      32'H3595: READ <= 8'H87;
      32'H3596: READ <= 8'H88;
      32'H3597: READ <= 8'H87;
      32'H3598: READ <= 8'H87;
      32'H3599: READ <= 8'H88;
      32'H3600: READ <= 8'H7b;
      32'H3601: READ <= 8'H7a;
      32'H3602: READ <= 8'H7b;
      32'H3603: READ <= 8'H7b;
      32'H3604: READ <= 8'H7b;
      32'H3605: READ <= 8'H7c;
      32'H3606: READ <= 8'H7d;
      32'H3607: READ <= 8'H7e;
      32'H3608: READ <= 8'H7f;
      32'H3609: READ <= 8'H7f;
      32'H3610: READ <= 8'H81;
      32'H3611: READ <= 8'H81;
      32'H3612: READ <= 8'H82;
      32'H3613: READ <= 8'H86;
      32'H3614: READ <= 8'H89;
      32'H3615: READ <= 8'H8d;
      32'H3616: READ <= 8'H91;
      32'H3617: READ <= 8'Ha1;
      32'H3618: READ <= 8'Hcc;
      32'H3619: READ <= 8'Hac;
      32'H3620: READ <= 8'H90;
      32'H3621: READ <= 8'H56;
      32'H3622: READ <= 8'H31;
      32'H3623: READ <= 8'H28;
      32'H3624: READ <= 8'H26;
      32'H3625: READ <= 8'H2d;
      32'H3626: READ <= 8'H28;
      32'H3627: READ <= 8'H22;
      32'H3628: READ <= 8'H21;
      32'H3629: READ <= 8'H25;
      32'H3630: READ <= 8'H27;
      32'H3631: READ <= 8'H1d;
      32'H3632: READ <= 8'H1c;
      32'H3633: READ <= 8'H21;
      32'H3634: READ <= 8'H18;
      32'H3635: READ <= 8'H65;
      32'H3636: READ <= 8'H6d;
      32'H3637: READ <= 8'H30;
      32'H3638: READ <= 8'H53;
      32'H3639: READ <= 8'H2a;
      32'H3640: READ <= 8'H8;
      32'H3641: READ <= 8'H8;
      32'H3642: READ <= 8'H46;
      32'H3643: READ <= 8'H71;
      32'H3644: READ <= 8'H36;
      32'H3645: READ <= 8'H3e;
      32'H3646: READ <= 8'H48;
      32'H3647: READ <= 8'H49;
      32'H3648: READ <= 8'H50;
      32'H3649: READ <= 8'H31;
      32'H3650: READ <= 8'H31;
      32'H3651: READ <= 8'H2f;
      32'H3652: READ <= 8'H53;
      32'H3653: READ <= 8'H4b;
      32'H3654: READ <= 8'Ha;
      32'H3655: READ <= 8'H6;
      32'H3656: READ <= 8'Ha;
      32'H3657: READ <= 8'H22;
      32'H3658: READ <= 8'H5d;
      32'H3659: READ <= 8'H7e;
      32'H3660: READ <= 8'H8c;
      32'H3661: READ <= 8'H9e;
      32'H3662: READ <= 8'H1d;
      32'H3663: READ <= 8'H2a;
      32'H3664: READ <= 8'H11;
      32'H3665: READ <= 8'H5f;
      32'H3666: READ <= 8'H7e;
      32'H3667: READ <= 8'H6d;
      32'H3668: READ <= 8'H6e;
      32'H3669: READ <= 8'H76;
      32'H3670: READ <= 8'H8a;
      32'H3671: READ <= 8'H93;
      32'H3672: READ <= 8'H96;
      32'H3673: READ <= 8'H95;
      32'H3674: READ <= 8'H95;
      32'H3675: READ <= 8'H92;
      32'H3676: READ <= 8'H71;
      32'H3677: READ <= 8'H7e;
      32'H3678: READ <= 8'H85;
      32'H3679: READ <= 8'H7e;
      32'H3680: READ <= 8'H7f;
      32'H3681: READ <= 8'H7f;
      32'H3682: READ <= 8'H80;
      32'H3683: READ <= 8'H81;
      32'H3684: READ <= 8'H81;
      32'H3685: READ <= 8'H82;
      32'H3686: READ <= 8'H86;
      32'H3687: READ <= 8'H71;
      32'H3688: READ <= 8'H8b;
      32'H3689: READ <= 8'H91;
      32'H3690: READ <= 8'H85;
      32'H3691: READ <= 8'H83;
      32'H3692: READ <= 8'H86;
      32'H3693: READ <= 8'H86;
      32'H3694: READ <= 8'H87;
      32'H3695: READ <= 8'H87;
      32'H3696: READ <= 8'H87;
      32'H3697: READ <= 8'H87;
      32'H3698: READ <= 8'H87;
      32'H3699: READ <= 8'H88;
      32'H3700: READ <= 8'H79;
      32'H3701: READ <= 8'H79;
      32'H3702: READ <= 8'H79;
      32'H3703: READ <= 8'H79;
      32'H3704: READ <= 8'H7a;
      32'H3705: READ <= 8'H7b;
      32'H3706: READ <= 8'H7c;
      32'H3707: READ <= 8'H7d;
      32'H3708: READ <= 8'H7e;
      32'H3709: READ <= 8'H7e;
      32'H3710: READ <= 8'H7f;
      32'H3711: READ <= 8'H80;
      32'H3712: READ <= 8'H80;
      32'H3713: READ <= 8'H83;
      32'H3714: READ <= 8'H85;
      32'H3715: READ <= 8'H88;
      32'H3716: READ <= 8'H90;
      32'H3717: READ <= 8'Hb1;
      32'H3718: READ <= 8'Hd1;
      32'H3719: READ <= 8'Hb2;
      32'H3720: READ <= 8'H89;
      32'H3721: READ <= 8'H71;
      32'H3722: READ <= 8'H4b;
      32'H3723: READ <= 8'H27;
      32'H3724: READ <= 8'H16;
      32'H3725: READ <= 8'H13;
      32'H3726: READ <= 8'H14;
      32'H3727: READ <= 8'H1c;
      32'H3728: READ <= 8'H28;
      32'H3729: READ <= 8'H30;
      32'H3730: READ <= 8'H49;
      32'H3731: READ <= 8'H5c;
      32'H3732: READ <= 8'H69;
      32'H3733: READ <= 8'H63;
      32'H3734: READ <= 8'H2b;
      32'H3735: READ <= 8'H6f;
      32'H3736: READ <= 8'H5e;
      32'H3737: READ <= 8'H29;
      32'H3738: READ <= 8'H4c;
      32'H3739: READ <= 8'H71;
      32'H3740: READ <= 8'H3c;
      32'H3741: READ <= 8'H11;
      32'H3742: READ <= 8'H15;
      32'H3743: READ <= 8'H5e;
      32'H3744: READ <= 8'H61;
      32'H3745: READ <= 8'H55;
      32'H3746: READ <= 8'H56;
      32'H3747: READ <= 8'H55;
      32'H3748: READ <= 8'H42;
      32'H3749: READ <= 8'H32;
      32'H3750: READ <= 8'H30;
      32'H3751: READ <= 8'H40;
      32'H3752: READ <= 8'H4e;
      32'H3753: READ <= 8'H41;
      32'H3754: READ <= 8'Hc;
      32'H3755: READ <= 8'H5;
      32'H3756: READ <= 8'H2;
      32'H3757: READ <= 8'H1d;
      32'H3758: READ <= 8'H4a;
      32'H3759: READ <= 8'H80;
      32'H3760: READ <= 8'H80;
      32'H3761: READ <= 8'H9d;
      32'H3762: READ <= 8'H4d;
      32'H3763: READ <= 8'H4d;
      32'H3764: READ <= 8'H1d;
      32'H3765: READ <= 8'H59;
      32'H3766: READ <= 8'H65;
      32'H3767: READ <= 8'H70;
      32'H3768: READ <= 8'H80;
      32'H3769: READ <= 8'H80;
      32'H3770: READ <= 8'H83;
      32'H3771: READ <= 8'H94;
      32'H3772: READ <= 8'H96;
      32'H3773: READ <= 8'H99;
      32'H3774: READ <= 8'H9d;
      32'H3775: READ <= 8'H89;
      32'H3776: READ <= 8'H85;
      32'H3777: READ <= 8'H82;
      32'H3778: READ <= 8'H8a;
      32'H3779: READ <= 8'H7f;
      32'H3780: READ <= 8'H7e;
      32'H3781: READ <= 8'H7e;
      32'H3782: READ <= 8'H7f;
      32'H3783: READ <= 8'H80;
      32'H3784: READ <= 8'H81;
      32'H3785: READ <= 8'H81;
      32'H3786: READ <= 8'H82;
      32'H3787: READ <= 8'H85;
      32'H3788: READ <= 8'H90;
      32'H3789: READ <= 8'Ha2;
      32'H3790: READ <= 8'H97;
      32'H3791: READ <= 8'H86;
      32'H3792: READ <= 8'H85;
      32'H3793: READ <= 8'H86;
      32'H3794: READ <= 8'H87;
      32'H3795: READ <= 8'H86;
      32'H3796: READ <= 8'H87;
      32'H3797: READ <= 8'H87;
      32'H3798: READ <= 8'H88;
      32'H3799: READ <= 8'H88;
      32'H3800: READ <= 8'H78;
      32'H3801: READ <= 8'H78;
      32'H3802: READ <= 8'H77;
      32'H3803: READ <= 8'H78;
      32'H3804: READ <= 8'H79;
      32'H3805: READ <= 8'H79;
      32'H3806: READ <= 8'H7b;
      32'H3807: READ <= 8'H7c;
      32'H3808: READ <= 8'H7c;
      32'H3809: READ <= 8'H7d;
      32'H3810: READ <= 8'H7d;
      32'H3811: READ <= 8'H7d;
      32'H3812: READ <= 8'H7f;
      32'H3813: READ <= 8'H80;
      32'H3814: READ <= 8'H82;
      32'H3815: READ <= 8'H84;
      32'H3816: READ <= 8'H89;
      32'H3817: READ <= 8'Ha2;
      32'H3818: READ <= 8'Hca;
      32'H3819: READ <= 8'Hb2;
      32'H3820: READ <= 8'H91;
      32'H3821: READ <= 8'H74;
      32'H3822: READ <= 8'H73;
      32'H3823: READ <= 8'H54;
      32'H3824: READ <= 8'H4d;
      32'H3825: READ <= 8'H43;
      32'H3826: READ <= 8'H44;
      32'H3827: READ <= 8'H4d;
      32'H3828: READ <= 8'H61;
      32'H3829: READ <= 8'H66;
      32'H3830: READ <= 8'H75;
      32'H3831: READ <= 8'H73;
      32'H3832: READ <= 8'H79;
      32'H3833: READ <= 8'H64;
      32'H3834: READ <= 8'H2e;
      32'H3835: READ <= 8'H5e;
      32'H3836: READ <= 8'H66;
      32'H3837: READ <= 8'H57;
      32'H3838: READ <= 8'H47;
      32'H3839: READ <= 8'H6c;
      32'H3840: READ <= 8'H7b;
      32'H3841: READ <= 8'H55;
      32'H3842: READ <= 8'H13;
      32'H3843: READ <= 8'H19;
      32'H3844: READ <= 8'H59;
      32'H3845: READ <= 8'H4f;
      32'H3846: READ <= 8'H42;
      32'H3847: READ <= 8'H4a;
      32'H3848: READ <= 8'H46;
      32'H3849: READ <= 8'H43;
      32'H3850: READ <= 8'H30;
      32'H3851: READ <= 8'H53;
      32'H3852: READ <= 8'H5d;
      32'H3853: READ <= 8'H24;
      32'H3854: READ <= 8'H19;
      32'H3855: READ <= 8'H20;
      32'H3856: READ <= 8'H7;
      32'H3857: READ <= 8'H23;
      32'H3858: READ <= 8'H43;
      32'H3859: READ <= 8'H7a;
      32'H3860: READ <= 8'H77;
      32'H3861: READ <= 8'H91;
      32'H3862: READ <= 8'H6f;
      32'H3863: READ <= 8'H68;
      32'H3864: READ <= 8'H2c;
      32'H3865: READ <= 8'H6f;
      32'H3866: READ <= 8'H5e;
      32'H3867: READ <= 8'H7a;
      32'H3868: READ <= 8'H8b;
      32'H3869: READ <= 8'H86;
      32'H3870: READ <= 8'H8b;
      32'H3871: READ <= 8'H8b;
      32'H3872: READ <= 8'H8a;
      32'H3873: READ <= 8'H9a;
      32'H3874: READ <= 8'Ha4;
      32'H3875: READ <= 8'H8f;
      32'H3876: READ <= 8'H81;
      32'H3877: READ <= 8'H98;
      32'H3878: READ <= 8'H8f;
      32'H3879: READ <= 8'H7e;
      32'H3880: READ <= 8'H7d;
      32'H3881: READ <= 8'H7e;
      32'H3882: READ <= 8'H7e;
      32'H3883: READ <= 8'H7f;
      32'H3884: READ <= 8'H80;
      32'H3885: READ <= 8'H81;
      32'H3886: READ <= 8'H82;
      32'H3887: READ <= 8'H82;
      32'H3888: READ <= 8'H8d;
      32'H3889: READ <= 8'H9a;
      32'H3890: READ <= 8'Ha6;
      32'H3891: READ <= 8'H99;
      32'H3892: READ <= 8'H8a;
      32'H3893: READ <= 8'H86;
      32'H3894: READ <= 8'H86;
      32'H3895: READ <= 8'H87;
      32'H3896: READ <= 8'H87;
      32'H3897: READ <= 8'H87;
      32'H3898: READ <= 8'H88;
      32'H3899: READ <= 8'H88;
      32'H3900: READ <= 8'H77;
      32'H3901: READ <= 8'H77;
      32'H3902: READ <= 8'H76;
      32'H3903: READ <= 8'H77;
      32'H3904: READ <= 8'H77;
      32'H3905: READ <= 8'H79;
      32'H3906: READ <= 8'H79;
      32'H3907: READ <= 8'H7a;
      32'H3908: READ <= 8'H7b;
      32'H3909: READ <= 8'H7b;
      32'H3910: READ <= 8'H7b;
      32'H3911: READ <= 8'H7d;
      32'H3912: READ <= 8'H7d;
      32'H3913: READ <= 8'H7e;
      32'H3914: READ <= 8'H7f;
      32'H3915: READ <= 8'H81;
      32'H3916: READ <= 8'H89;
      32'H3917: READ <= 8'Haf;
      32'H3918: READ <= 8'Hcf;
      32'H3919: READ <= 8'Hb6;
      32'H3920: READ <= 8'H7c;
      32'H3921: READ <= 8'H86;
      32'H3922: READ <= 8'H6a;
      32'H3923: READ <= 8'H6b;
      32'H3924: READ <= 8'H59;
      32'H3925: READ <= 8'H4e;
      32'H3926: READ <= 8'H4d;
      32'H3927: READ <= 8'H51;
      32'H3928: READ <= 8'H62;
      32'H3929: READ <= 8'H76;
      32'H3930: READ <= 8'H70;
      32'H3931: READ <= 8'H71;
      32'H3932: READ <= 8'H7d;
      32'H3933: READ <= 8'H72;
      32'H3934: READ <= 8'H37;
      32'H3935: READ <= 8'H64;
      32'H3936: READ <= 8'H6b;
      32'H3937: READ <= 8'H6a;
      32'H3938: READ <= 8'H35;
      32'H3939: READ <= 8'H4a;
      32'H3940: READ <= 8'H77;
      32'H3941: READ <= 8'H77;
      32'H3942: READ <= 8'H4c;
      32'H3943: READ <= 8'H15;
      32'H3944: READ <= 8'H15;
      32'H3945: READ <= 8'H49;
      32'H3946: READ <= 8'H6c;
      32'H3947: READ <= 8'H3a;
      32'H3948: READ <= 8'H35;
      32'H3949: READ <= 8'H4b;
      32'H3950: READ <= 8'H2e;
      32'H3951: READ <= 8'H46;
      32'H3952: READ <= 8'H6b;
      32'H3953: READ <= 8'H8;
      32'H3954: READ <= 8'H51;
      32'H3955: READ <= 8'H94;
      32'H3956: READ <= 8'H48;
      32'H3957: READ <= 8'H33;
      32'H3958: READ <= 8'H36;
      32'H3959: READ <= 8'H70;
      32'H3960: READ <= 8'H70;
      32'H3961: READ <= 8'H92;
      32'H3962: READ <= 8'H72;
      32'H3963: READ <= 8'H6d;
      32'H3964: READ <= 8'H33;
      32'H3965: READ <= 8'H5d;
      32'H3966: READ <= 8'H46;
      32'H3967: READ <= 8'H6a;
      32'H3968: READ <= 8'H8e;
      32'H3969: READ <= 8'H7f;
      32'H3970: READ <= 8'H81;
      32'H3971: READ <= 8'H83;
      32'H3972: READ <= 8'H8e;
      32'H3973: READ <= 8'H92;
      32'H3974: READ <= 8'H99;
      32'H3975: READ <= 8'H94;
      32'H3976: READ <= 8'H88;
      32'H3977: READ <= 8'Ha5;
      32'H3978: READ <= 8'H97;
      32'H3979: READ <= 8'H7f;
      32'H3980: READ <= 8'H7d;
      32'H3981: READ <= 8'H7d;
      32'H3982: READ <= 8'H7d;
      32'H3983: READ <= 8'H7f;
      32'H3984: READ <= 8'H7f;
      32'H3985: READ <= 8'H80;
      32'H3986: READ <= 8'H82;
      32'H3987: READ <= 8'H82;
      32'H3988: READ <= 8'H84;
      32'H3989: READ <= 8'H92;
      32'H3990: READ <= 8'Ha1;
      32'H3991: READ <= 8'Ha8;
      32'H3992: READ <= 8'Ha0;
      32'H3993: READ <= 8'H8d;
      32'H3994: READ <= 8'H86;
      32'H3995: READ <= 8'H88;
      32'H3996: READ <= 8'H87;
      32'H3997: READ <= 8'H87;
      32'H3998: READ <= 8'H88;
      32'H3999: READ <= 8'H88;
      32'H4000: READ <= 8'H76;
      32'H4001: READ <= 8'H76;
      32'H4002: READ <= 8'H75;
      32'H4003: READ <= 8'H76;
      32'H4004: READ <= 8'H76;
      32'H4005: READ <= 8'H77;
      32'H4006: READ <= 8'H77;
      32'H4007: READ <= 8'H78;
      32'H4008: READ <= 8'H79;
      32'H4009: READ <= 8'H7a;
      32'H4010: READ <= 8'H7a;
      32'H4011: READ <= 8'H7b;
      32'H4012: READ <= 8'H7c;
      32'H4013: READ <= 8'H7c;
      32'H4014: READ <= 8'H7c;
      32'H4015: READ <= 8'H7f;
      32'H4016: READ <= 8'H85;
      32'H4017: READ <= 8'Ha9;
      32'H4018: READ <= 8'Hc8;
      32'H4019: READ <= 8'Hb0;
      32'H4020: READ <= 8'H8c;
      32'H4021: READ <= 8'H75;
      32'H4022: READ <= 8'H69;
      32'H4023: READ <= 8'H6e;
      32'H4024: READ <= 8'H48;
      32'H4025: READ <= 8'H4b;
      32'H4026: READ <= 8'H4c;
      32'H4027: READ <= 8'H5c;
      32'H4028: READ <= 8'H5a;
      32'H4029: READ <= 8'H6d;
      32'H4030: READ <= 8'H60;
      32'H4031: READ <= 8'H57;
      32'H4032: READ <= 8'H60;
      32'H4033: READ <= 8'H64;
      32'H4034: READ <= 8'H3e;
      32'H4035: READ <= 8'H61;
      32'H4036: READ <= 8'H65;
      32'H4037: READ <= 8'H6f;
      32'H4038: READ <= 8'H48;
      32'H4039: READ <= 8'H24;
      32'H4040: READ <= 8'H60;
      32'H4041: READ <= 8'H69;
      32'H4042: READ <= 8'H65;
      32'H4043: READ <= 8'H53;
      32'H4044: READ <= 8'H2a;
      32'H4045: READ <= 8'H1a;
      32'H4046: READ <= 8'H42;
      32'H4047: READ <= 8'H1c;
      32'H4048: READ <= 8'H18;
      32'H4049: READ <= 8'H34;
      32'H4050: READ <= 8'H2a;
      32'H4051: READ <= 8'H37;
      32'H4052: READ <= 8'H5b;
      32'H4053: READ <= 8'H3;
      32'H4054: READ <= 8'H95;
      32'H4055: READ <= 8'Hb7;
      32'H4056: READ <= 8'Ha3;
      32'H4057: READ <= 8'H6f;
      32'H4058: READ <= 8'H41;
      32'H4059: READ <= 8'H65;
      32'H4060: READ <= 8'H70;
      32'H4061: READ <= 8'H95;
      32'H4062: READ <= 8'H5d;
      32'H4063: READ <= 8'H5f;
      32'H4064: READ <= 8'H46;
      32'H4065: READ <= 8'H61;
      32'H4066: READ <= 8'H5b;
      32'H4067: READ <= 8'H5c;
      32'H4068: READ <= 8'H7c;
      32'H4069: READ <= 8'H81;
      32'H4070: READ <= 8'H82;
      32'H4071: READ <= 8'H89;
      32'H4072: READ <= 8'H8d;
      32'H4073: READ <= 8'H95;
      32'H4074: READ <= 8'H96;
      32'H4075: READ <= 8'H93;
      32'H4076: READ <= 8'H93;
      32'H4077: READ <= 8'Ha2;
      32'H4078: READ <= 8'H94;
      32'H4079: READ <= 8'H7f;
      32'H4080: READ <= 8'H7c;
      32'H4081: READ <= 8'H7c;
      32'H4082: READ <= 8'H7d;
      32'H4083: READ <= 8'H7e;
      32'H4084: READ <= 8'H7f;
      32'H4085: READ <= 8'H80;
      32'H4086: READ <= 8'H81;
      32'H4087: READ <= 8'H82;
      32'H4088: READ <= 8'H82;
      32'H4089: READ <= 8'H88;
      32'H4090: READ <= 8'H9f;
      32'H4091: READ <= 8'Ha5;
      32'H4092: READ <= 8'Haf;
      32'H4093: READ <= 8'Ha9;
      32'H4094: READ <= 8'H93;
      32'H4095: READ <= 8'H88;
      32'H4096: READ <= 8'H88;
      32'H4097: READ <= 8'H88;
      32'H4098: READ <= 8'H88;
      32'H4099: READ <= 8'H88;
      32'H4100: READ <= 8'H75;
      32'H4101: READ <= 8'H75;
      32'H4102: READ <= 8'H74;
      32'H4103: READ <= 8'H75;
      32'H4104: READ <= 8'H75;
      32'H4105: READ <= 8'H76;
      32'H4106: READ <= 8'H77;
      32'H4107: READ <= 8'H76;
      32'H4108: READ <= 8'H77;
      32'H4109: READ <= 8'H78;
      32'H4110: READ <= 8'H79;
      32'H4111: READ <= 8'H79;
      32'H4112: READ <= 8'H7a;
      32'H4113: READ <= 8'H7a;
      32'H4114: READ <= 8'H7c;
      32'H4115: READ <= 8'H7c;
      32'H4116: READ <= 8'H81;
      32'H4117: READ <= 8'H9a;
      32'H4118: READ <= 8'Hbc;
      32'H4119: READ <= 8'Ha8;
      32'H4120: READ <= 8'H8c;
      32'H4121: READ <= 8'H7d;
      32'H4122: READ <= 8'H68;
      32'H4123: READ <= 8'H62;
      32'H4124: READ <= 8'H58;
      32'H4125: READ <= 8'H53;
      32'H4126: READ <= 8'H4e;
      32'H4127: READ <= 8'H63;
      32'H4128: READ <= 8'H5d;
      32'H4129: READ <= 8'H5e;
      32'H4130: READ <= 8'H68;
      32'H4131: READ <= 8'H5e;
      32'H4132: READ <= 8'H74;
      32'H4133: READ <= 8'H69;
      32'H4134: READ <= 8'H55;
      32'H4135: READ <= 8'H42;
      32'H4136: READ <= 8'H5c;
      32'H4137: READ <= 8'H61;
      32'H4138: READ <= 8'H60;
      32'H4139: READ <= 8'H1e;
      32'H4140: READ <= 8'H3a;
      32'H4141: READ <= 8'H59;
      32'H4142: READ <= 8'H53;
      32'H4143: READ <= 8'H62;
      32'H4144: READ <= 8'H5e;
      32'H4145: READ <= 8'H1b;
      32'H4146: READ <= 8'He;
      32'H4147: READ <= 8'H3;
      32'H4148: READ <= 8'H6;
      32'H4149: READ <= 8'H23;
      32'H4150: READ <= 8'H21;
      32'H4151: READ <= 8'H1e;
      32'H4152: READ <= 8'H2c;
      32'H4153: READ <= 8'H51;
      32'H4154: READ <= 8'Hdb;
      32'H4155: READ <= 8'Ha9;
      32'H4156: READ <= 8'H8a;
      32'H4157: READ <= 8'H8a;
      32'H4158: READ <= 8'H44;
      32'H4159: READ <= 8'H60;
      32'H4160: READ <= 8'H6c;
      32'H4161: READ <= 8'H90;
      32'H4162: READ <= 8'H49;
      32'H4163: READ <= 8'H4c;
      32'H4164: READ <= 8'H49;
      32'H4165: READ <= 8'H69;
      32'H4166: READ <= 8'H71;
      32'H4167: READ <= 8'H66;
      32'H4168: READ <= 8'H77;
      32'H4169: READ <= 8'H76;
      32'H4170: READ <= 8'H7b;
      32'H4171: READ <= 8'H81;
      32'H4172: READ <= 8'H85;
      32'H4173: READ <= 8'H91;
      32'H4174: READ <= 8'H9b;
      32'H4175: READ <= 8'H99;
      32'H4176: READ <= 8'Ha1;
      32'H4177: READ <= 8'Ha8;
      32'H4178: READ <= 8'H97;
      32'H4179: READ <= 8'H7e;
      32'H4180: READ <= 8'H7c;
      32'H4181: READ <= 8'H7c;
      32'H4182: READ <= 8'H7d;
      32'H4183: READ <= 8'H7e;
      32'H4184: READ <= 8'H7f;
      32'H4185: READ <= 8'H7f;
      32'H4186: READ <= 8'H80;
      32'H4187: READ <= 8'H82;
      32'H4188: READ <= 8'H82;
      32'H4189: READ <= 8'H83;
      32'H4190: READ <= 8'H8f;
      32'H4191: READ <= 8'H9c;
      32'H4192: READ <= 8'H96;
      32'H4193: READ <= 8'Ha3;
      32'H4194: READ <= 8'H95;
      32'H4195: READ <= 8'H88;
      32'H4196: READ <= 8'H88;
      32'H4197: READ <= 8'H89;
      32'H4198: READ <= 8'H88;
      32'H4199: READ <= 8'H89;
      32'H4200: READ <= 8'H74;
      32'H4201: READ <= 8'H74;
      32'H4202: READ <= 8'H74;
      32'H4203: READ <= 8'H75;
      32'H4204: READ <= 8'H74;
      32'H4205: READ <= 8'H76;
      32'H4206: READ <= 8'H76;
      32'H4207: READ <= 8'H75;
      32'H4208: READ <= 8'H76;
      32'H4209: READ <= 8'H76;
      32'H4210: READ <= 8'H77;
      32'H4211: READ <= 8'H78;
      32'H4212: READ <= 8'H78;
      32'H4213: READ <= 8'H79;
      32'H4214: READ <= 8'H7a;
      32'H4215: READ <= 8'H7b;
      32'H4216: READ <= 8'H7d;
      32'H4217: READ <= 8'H95;
      32'H4218: READ <= 8'Hbc;
      32'H4219: READ <= 8'Hb0;
      32'H4220: READ <= 8'H89;
      32'H4221: READ <= 8'H6f;
      32'H4222: READ <= 8'H7a;
      32'H4223: READ <= 8'H6f;
      32'H4224: READ <= 8'H4e;
      32'H4225: READ <= 8'H48;
      32'H4226: READ <= 8'H3f;
      32'H4227: READ <= 8'H52;
      32'H4228: READ <= 8'H56;
      32'H4229: READ <= 8'H4d;
      32'H4230: READ <= 8'H4d;
      32'H4231: READ <= 8'H57;
      32'H4232: READ <= 8'H60;
      32'H4233: READ <= 8'H4f;
      32'H4234: READ <= 8'H3c;
      32'H4235: READ <= 8'H32;
      32'H4236: READ <= 8'H55;
      32'H4237: READ <= 8'H56;
      32'H4238: READ <= 8'H64;
      32'H4239: READ <= 8'H1a;
      32'H4240: READ <= 8'H1d;
      32'H4241: READ <= 8'H4e;
      32'H4242: READ <= 8'H59;
      32'H4243: READ <= 8'H47;
      32'H4244: READ <= 8'H42;
      32'H4245: READ <= 8'H23;
      32'H4246: READ <= 8'H18;
      32'H4247: READ <= 8'H8;
      32'H4248: READ <= 8'H11;
      32'H4249: READ <= 8'H31;
      32'H4250: READ <= 8'H33;
      32'H4251: READ <= 8'H9;
      32'H4252: READ <= 8'H1e;
      32'H4253: READ <= 8'Hcd;
      32'H4254: READ <= 8'Hfc;
      32'H4255: READ <= 8'Ha4;
      32'H4256: READ <= 8'H66;
      32'H4257: READ <= 8'H76;
      32'H4258: READ <= 8'H3a;
      32'H4259: READ <= 8'H5b;
      32'H4260: READ <= 8'H69;
      32'H4261: READ <= 8'H7e;
      32'H4262: READ <= 8'H30;
      32'H4263: READ <= 8'H3d;
      32'H4264: READ <= 8'H47;
      32'H4265: READ <= 8'H5d;
      32'H4266: READ <= 8'H68;
      32'H4267: READ <= 8'H6b;
      32'H4268: READ <= 8'H6c;
      32'H4269: READ <= 8'H69;
      32'H4270: READ <= 8'H6f;
      32'H4271: READ <= 8'H6c;
      32'H4272: READ <= 8'H88;
      32'H4273: READ <= 8'H8e;
      32'H4274: READ <= 8'H9d;
      32'H4275: READ <= 8'Ha9;
      32'H4276: READ <= 8'Ha4;
      32'H4277: READ <= 8'Ha8;
      32'H4278: READ <= 8'H9e;
      32'H4279: READ <= 8'H80;
      32'H4280: READ <= 8'H7b;
      32'H4281: READ <= 8'H7c;
      32'H4282: READ <= 8'H7c;
      32'H4283: READ <= 8'H7d;
      32'H4284: READ <= 8'H7e;
      32'H4285: READ <= 8'H7f;
      32'H4286: READ <= 8'H81;
      32'H4287: READ <= 8'H82;
      32'H4288: READ <= 8'H82;
      32'H4289: READ <= 8'H83;
      32'H4290: READ <= 8'H83;
      32'H4291: READ <= 8'H8a;
      32'H4292: READ <= 8'H86;
      32'H4293: READ <= 8'H8a;
      32'H4294: READ <= 8'H89;
      32'H4295: READ <= 8'H88;
      32'H4296: READ <= 8'H88;
      32'H4297: READ <= 8'H88;
      32'H4298: READ <= 8'H89;
      32'H4299: READ <= 8'H89;
      32'H4300: READ <= 8'H74;
      32'H4301: READ <= 8'H73;
      32'H4302: READ <= 8'H73;
      32'H4303: READ <= 8'H74;
      32'H4304: READ <= 8'H74;
      32'H4305: READ <= 8'H75;
      32'H4306: READ <= 8'H75;
      32'H4307: READ <= 8'H75;
      32'H4308: READ <= 8'H74;
      32'H4309: READ <= 8'H75;
      32'H4310: READ <= 8'H75;
      32'H4311: READ <= 8'H76;
      32'H4312: READ <= 8'H76;
      32'H4313: READ <= 8'H77;
      32'H4314: READ <= 8'H78;
      32'H4315: READ <= 8'H79;
      32'H4316: READ <= 8'H81;
      32'H4317: READ <= 8'H9e;
      32'H4318: READ <= 8'Hc3;
      32'H4319: READ <= 8'Hbd;
      32'H4320: READ <= 8'H89;
      32'H4321: READ <= 8'H51;
      32'H4322: READ <= 8'H79;
      32'H4323: READ <= 8'H6f;
      32'H4324: READ <= 8'H53;
      32'H4325: READ <= 8'H46;
      32'H4326: READ <= 8'H35;
      32'H4327: READ <= 8'H36;
      32'H4328: READ <= 8'H30;
      32'H4329: READ <= 8'H2e;
      32'H4330: READ <= 8'H30;
      32'H4331: READ <= 8'H34;
      32'H4332: READ <= 8'H2e;
      32'H4333: READ <= 8'H38;
      32'H4334: READ <= 8'H35;
      32'H4335: READ <= 8'H2b;
      32'H4336: READ <= 8'H4a;
      32'H4337: READ <= 8'H56;
      32'H4338: READ <= 8'H50;
      32'H4339: READ <= 8'H2a;
      32'H4340: READ <= 8'H10;
      32'H4341: READ <= 8'H37;
      32'H4342: READ <= 8'H52;
      32'H4343: READ <= 8'H36;
      32'H4344: READ <= 8'H1e;
      32'H4345: READ <= 8'H17;
      32'H4346: READ <= 8'H1a;
      32'H4347: READ <= 8'Hf;
      32'H4348: READ <= 8'H40;
      32'H4349: READ <= 8'H50;
      32'H4350: READ <= 8'H36;
      32'H4351: READ <= 8'H1;
      32'H4352: READ <= 8'H2a;
      32'H4353: READ <= 8'He6;
      32'H4354: READ <= 8'Hf7;
      32'H4355: READ <= 8'Hb5;
      32'H4356: READ <= 8'H5b;
      32'H4357: READ <= 8'H75;
      32'H4358: READ <= 8'H36;
      32'H4359: READ <= 8'H51;
      32'H4360: READ <= 8'H6c;
      32'H4361: READ <= 8'H76;
      32'H4362: READ <= 8'H1c;
      32'H4363: READ <= 8'H36;
      32'H4364: READ <= 8'H4a;
      32'H4365: READ <= 8'H5c;
      32'H4366: READ <= 8'H68;
      32'H4367: READ <= 8'H67;
      32'H4368: READ <= 8'H72;
      32'H4369: READ <= 8'H6e;
      32'H4370: READ <= 8'H69;
      32'H4371: READ <= 8'H69;
      32'H4372: READ <= 8'H84;
      32'H4373: READ <= 8'H90;
      32'H4374: READ <= 8'H98;
      32'H4375: READ <= 8'H97;
      32'H4376: READ <= 8'Ha7;
      32'H4377: READ <= 8'Hb3;
      32'H4378: READ <= 8'H9c;
      32'H4379: READ <= 8'H7f;
      32'H4380: READ <= 8'H7c;
      32'H4381: READ <= 8'H7b;
      32'H4382: READ <= 8'H7d;
      32'H4383: READ <= 8'H7d;
      32'H4384: READ <= 8'H7e;
      32'H4385: READ <= 8'H7f;
      32'H4386: READ <= 8'H81;
      32'H4387: READ <= 8'H81;
      32'H4388: READ <= 8'H82;
      32'H4389: READ <= 8'H83;
      32'H4390: READ <= 8'H84;
      32'H4391: READ <= 8'H85;
      32'H4392: READ <= 8'H86;
      32'H4393: READ <= 8'H87;
      32'H4394: READ <= 8'H88;
      32'H4395: READ <= 8'H88;
      32'H4396: READ <= 8'H88;
      32'H4397: READ <= 8'H89;
      32'H4398: READ <= 8'H89;
      32'H4399: READ <= 8'H88;
      32'H4400: READ <= 8'H73;
      32'H4401: READ <= 8'H73;
      32'H4402: READ <= 8'H73;
      32'H4403: READ <= 8'H73;
      32'H4404: READ <= 8'H73;
      32'H4405: READ <= 8'H74;
      32'H4406: READ <= 8'H75;
      32'H4407: READ <= 8'H75;
      32'H4408: READ <= 8'H74;
      32'H4409: READ <= 8'H74;
      32'H4410: READ <= 8'H74;
      32'H4411: READ <= 8'H75;
      32'H4412: READ <= 8'H75;
      32'H4413: READ <= 8'H76;
      32'H4414: READ <= 8'H77;
      32'H4415: READ <= 8'H78;
      32'H4416: READ <= 8'H7c;
      32'H4417: READ <= 8'H8e;
      32'H4418: READ <= 8'Hcb;
      32'H4419: READ <= 8'Hc7;
      32'H4420: READ <= 8'H91;
      32'H4421: READ <= 8'H57;
      32'H4422: READ <= 8'H6a;
      32'H4423: READ <= 8'H63;
      32'H4424: READ <= 8'H61;
      32'H4425: READ <= 8'H37;
      32'H4426: READ <= 8'H3f;
      32'H4427: READ <= 8'H3d;
      32'H4428: READ <= 8'H39;
      32'H4429: READ <= 8'H34;
      32'H4430: READ <= 8'H34;
      32'H4431: READ <= 8'H41;
      32'H4432: READ <= 8'H44;
      32'H4433: READ <= 8'H34;
      32'H4434: READ <= 8'H20;
      32'H4435: READ <= 8'H16;
      32'H4436: READ <= 8'H48;
      32'H4437: READ <= 8'H54;
      32'H4438: READ <= 8'H44;
      32'H4439: READ <= 8'H47;
      32'H4440: READ <= 8'H8;
      32'H4441: READ <= 8'H26;
      32'H4442: READ <= 8'H42;
      32'H4443: READ <= 8'H2d;
      32'H4444: READ <= 8'H18;
      32'H4445: READ <= 8'He;
      32'H4446: READ <= 8'H19;
      32'H4447: READ <= 8'H42;
      32'H4448: READ <= 8'H48;
      32'H4449: READ <= 8'H71;
      32'H4450: READ <= 8'H21;
      32'H4451: READ <= 8'H23;
      32'H4452: READ <= 8'H9e;
      32'H4453: READ <= 8'Hda;
      32'H4454: READ <= 8'He6;
      32'H4455: READ <= 8'Hca;
      32'H4456: READ <= 8'H6c;
      32'H4457: READ <= 8'H5f;
      32'H4458: READ <= 8'H2a;
      32'H4459: READ <= 8'H4f;
      32'H4460: READ <= 8'H6b;
      32'H4461: READ <= 8'H7c;
      32'H4462: READ <= 8'H24;
      32'H4463: READ <= 8'H2f;
      32'H4464: READ <= 8'H41;
      32'H4465: READ <= 8'H5b;
      32'H4466: READ <= 8'H62;
      32'H4467: READ <= 8'H65;
      32'H4468: READ <= 8'H65;
      32'H4469: READ <= 8'H62;
      32'H4470: READ <= 8'H75;
      32'H4471: READ <= 8'H71;
      32'H4472: READ <= 8'H90;
      32'H4473: READ <= 8'H94;
      32'H4474: READ <= 8'H9d;
      32'H4475: READ <= 8'Ha6;
      32'H4476: READ <= 8'Ha2;
      32'H4477: READ <= 8'Hb0;
      32'H4478: READ <= 8'H96;
      32'H4479: READ <= 8'H7e;
      32'H4480: READ <= 8'H7b;
      32'H4481: READ <= 8'H7b;
      32'H4482: READ <= 8'H7d;
      32'H4483: READ <= 8'H7e;
      32'H4484: READ <= 8'H7e;
      32'H4485: READ <= 8'H7f;
      32'H4486: READ <= 8'H81;
      32'H4487: READ <= 8'H81;
      32'H4488: READ <= 8'H82;
      32'H4489: READ <= 8'H83;
      32'H4490: READ <= 8'H84;
      32'H4491: READ <= 8'H85;
      32'H4492: READ <= 8'H86;
      32'H4493: READ <= 8'H86;
      32'H4494: READ <= 8'H88;
      32'H4495: READ <= 8'H88;
      32'H4496: READ <= 8'H88;
      32'H4497: READ <= 8'H89;
      32'H4498: READ <= 8'H89;
      32'H4499: READ <= 8'H89;
      32'H4500: READ <= 8'H73;
      32'H4501: READ <= 8'H72;
      32'H4502: READ <= 8'H72;
      32'H4503: READ <= 8'H73;
      32'H4504: READ <= 8'H73;
      32'H4505: READ <= 8'H74;
      32'H4506: READ <= 8'H75;
      32'H4507: READ <= 8'H74;
      32'H4508: READ <= 8'H74;
      32'H4509: READ <= 8'H74;
      32'H4510: READ <= 8'H74;
      32'H4511: READ <= 8'H74;
      32'H4512: READ <= 8'H74;
      32'H4513: READ <= 8'H75;
      32'H4514: READ <= 8'H76;
      32'H4515: READ <= 8'H78;
      32'H4516: READ <= 8'H80;
      32'H4517: READ <= 8'H9e;
      32'H4518: READ <= 8'Hbd;
      32'H4519: READ <= 8'Hb8;
      32'H4520: READ <= 8'Hae;
      32'H4521: READ <= 8'H83;
      32'H4522: READ <= 8'H78;
      32'H4523: READ <= 8'H6b;
      32'H4524: READ <= 8'H57;
      32'H4525: READ <= 8'H4a;
      32'H4526: READ <= 8'H48;
      32'H4527: READ <= 8'H3a;
      32'H4528: READ <= 8'H30;
      32'H4529: READ <= 8'H24;
      32'H4530: READ <= 8'H1c;
      32'H4531: READ <= 8'H1a;
      32'H4532: READ <= 8'H26;
      32'H4533: READ <= 8'H2f;
      32'H4534: READ <= 8'H2d;
      32'H4535: READ <= 8'Hc;
      32'H4536: READ <= 8'H37;
      32'H4537: READ <= 8'H48;
      32'H4538: READ <= 8'H33;
      32'H4539: READ <= 8'H4c;
      32'H4540: READ <= 8'Hc;
      32'H4541: READ <= 8'H16;
      32'H4542: READ <= 8'H2e;
      32'H4543: READ <= 8'H34;
      32'H4544: READ <= 8'H1e;
      32'H4545: READ <= 8'H26;
      32'H4546: READ <= 8'H6f;
      32'H4547: READ <= 8'Ha1;
      32'H4548: READ <= 8'Ha0;
      32'H4549: READ <= 8'H8d;
      32'H4550: READ <= 8'H4d;
      32'H4551: READ <= 8'H68;
      32'H4552: READ <= 8'Ha5;
      32'H4553: READ <= 8'Hc9;
      32'H4554: READ <= 8'Hd1;
      32'H4555: READ <= 8'Hca;
      32'H4556: READ <= 8'H78;
      32'H4557: READ <= 8'H4f;
      32'H4558: READ <= 8'H18;
      32'H4559: READ <= 8'H46;
      32'H4560: READ <= 8'H6b;
      32'H4561: READ <= 8'H88;
      32'H4562: READ <= 8'H43;
      32'H4563: READ <= 8'H36;
      32'H4564: READ <= 8'H4c;
      32'H4565: READ <= 8'H59;
      32'H4566: READ <= 8'H5e;
      32'H4567: READ <= 8'H6f;
      32'H4568: READ <= 8'H62;
      32'H4569: READ <= 8'H6e;
      32'H4570: READ <= 8'H72;
      32'H4571: READ <= 8'H71;
      32'H4572: READ <= 8'H7f;
      32'H4573: READ <= 8'H8a;
      32'H4574: READ <= 8'H92;
      32'H4575: READ <= 8'H9a;
      32'H4576: READ <= 8'Hac;
      32'H4577: READ <= 8'Had;
      32'H4578: READ <= 8'H93;
      32'H4579: READ <= 8'H7d;
      32'H4580: READ <= 8'H7b;
      32'H4581: READ <= 8'H7b;
      32'H4582: READ <= 8'H7c;
      32'H4583: READ <= 8'H7d;
      32'H4584: READ <= 8'H7e;
      32'H4585: READ <= 8'H7f;
      32'H4586: READ <= 8'H81;
      32'H4587: READ <= 8'H82;
      32'H4588: READ <= 8'H82;
      32'H4589: READ <= 8'H83;
      32'H4590: READ <= 8'H84;
      32'H4591: READ <= 8'H85;
      32'H4592: READ <= 8'H86;
      32'H4593: READ <= 8'H86;
      32'H4594: READ <= 8'H88;
      32'H4595: READ <= 8'H89;
      32'H4596: READ <= 8'H89;
      32'H4597: READ <= 8'H89;
      32'H4598: READ <= 8'H89;
      32'H4599: READ <= 8'H89;
      32'H4600: READ <= 8'H72;
      32'H4601: READ <= 8'H72;
      32'H4602: READ <= 8'H71;
      32'H4603: READ <= 8'H72;
      32'H4604: READ <= 8'H72;
      32'H4605: READ <= 8'H73;
      32'H4606: READ <= 8'H74;
      32'H4607: READ <= 8'H74;
      32'H4608: READ <= 8'H73;
      32'H4609: READ <= 8'H73;
      32'H4610: READ <= 8'H73;
      32'H4611: READ <= 8'H74;
      32'H4612: READ <= 8'H74;
      32'H4613: READ <= 8'H74;
      32'H4614: READ <= 8'H76;
      32'H4615: READ <= 8'H77;
      32'H4616: READ <= 8'H7a;
      32'H4617: READ <= 8'H89;
      32'H4618: READ <= 8'H9f;
      32'H4619: READ <= 8'Ha0;
      32'H4620: READ <= 8'Hb1;
      32'H4621: READ <= 8'H90;
      32'H4622: READ <= 8'H86;
      32'H4623: READ <= 8'H6c;
      32'H4624: READ <= 8'H51;
      32'H4625: READ <= 8'H54;
      32'H4626: READ <= 8'H47;
      32'H4627: READ <= 8'H35;
      32'H4628: READ <= 8'H2c;
      32'H4629: READ <= 8'H22;
      32'H4630: READ <= 8'H1a;
      32'H4631: READ <= 8'H16;
      32'H4632: READ <= 8'H15;
      32'H4633: READ <= 8'H15;
      32'H4634: READ <= 8'H14;
      32'H4635: READ <= 8'Hb;
      32'H4636: READ <= 8'H27;
      32'H4637: READ <= 8'H43;
      32'H4638: READ <= 8'H1c;
      32'H4639: READ <= 8'H50;
      32'H4640: READ <= 8'He;
      32'H4641: READ <= 8'Hd;
      32'H4642: READ <= 8'H17;
      32'H4643: READ <= 8'H30;
      32'H4644: READ <= 8'H5f;
      32'H4645: READ <= 8'Hc3;
      32'H4646: READ <= 8'Hef;
      32'H4647: READ <= 8'Hf1;
      32'H4648: READ <= 8'Hda;
      32'H4649: READ <= 8'Hb7;
      32'H4650: READ <= 8'Haf;
      32'H4651: READ <= 8'H9a;
      32'H4652: READ <= 8'Ha1;
      32'H4653: READ <= 8'Hb3;
      32'H4654: READ <= 8'Hb4;
      32'H4655: READ <= 8'Hbe;
      32'H4656: READ <= 8'H82;
      32'H4657: READ <= 8'H59;
      32'H4658: READ <= 8'H2f;
      32'H4659: READ <= 8'H26;
      32'H4660: READ <= 8'H54;
      32'H4661: READ <= 8'H8f;
      32'H4662: READ <= 8'H61;
      32'H4663: READ <= 8'H5d;
      32'H4664: READ <= 8'H3c;
      32'H4665: READ <= 8'H56;
      32'H4666: READ <= 8'H6d;
      32'H4667: READ <= 8'H6c;
      32'H4668: READ <= 8'H7f;
      32'H4669: READ <= 8'H71;
      32'H4670: READ <= 8'H7e;
      32'H4671: READ <= 8'H85;
      32'H4672: READ <= 8'H8b;
      32'H4673: READ <= 8'H92;
      32'H4674: READ <= 8'H9c;
      32'H4675: READ <= 8'Ha1;
      32'H4676: READ <= 8'H9f;
      32'H4677: READ <= 8'Ha9;
      32'H4678: READ <= 8'H8c;
      32'H4679: READ <= 8'H7b;
      32'H4680: READ <= 8'H7a;
      32'H4681: READ <= 8'H7b;
      32'H4682: READ <= 8'H7c;
      32'H4683: READ <= 8'H7d;
      32'H4684: READ <= 8'H7d;
      32'H4685: READ <= 8'H7f;
      32'H4686: READ <= 8'H80;
      32'H4687: READ <= 8'H81;
      32'H4688: READ <= 8'H82;
      32'H4689: READ <= 8'H83;
      32'H4690: READ <= 8'H84;
      32'H4691: READ <= 8'H85;
      32'H4692: READ <= 8'H86;
      32'H4693: READ <= 8'H87;
      32'H4694: READ <= 8'H89;
      32'H4695: READ <= 8'H89;
      32'H4696: READ <= 8'H89;
      32'H4697: READ <= 8'H89;
      32'H4698: READ <= 8'H8a;
      32'H4699: READ <= 8'H8a;
      32'H4700: READ <= 8'H71;
      32'H4701: READ <= 8'H71;
      32'H4702: READ <= 8'H71;
      32'H4703: READ <= 8'H71;
      32'H4704: READ <= 8'H72;
      32'H4705: READ <= 8'H72;
      32'H4706: READ <= 8'H73;
      32'H4707: READ <= 8'H73;
      32'H4708: READ <= 8'H73;
      32'H4709: READ <= 8'H73;
      32'H4710: READ <= 8'H73;
      32'H4711: READ <= 8'H73;
      32'H4712: READ <= 8'H73;
      32'H4713: READ <= 8'H74;
      32'H4714: READ <= 8'H74;
      32'H4715: READ <= 8'H75;
      32'H4716: READ <= 8'H78;
      32'H4717: READ <= 8'H82;
      32'H4718: READ <= 8'H85;
      32'H4719: READ <= 8'Ha6;
      32'H4720: READ <= 8'Hb9;
      32'H4721: READ <= 8'Hc3;
      32'H4722: READ <= 8'Ha5;
      32'H4723: READ <= 8'H83;
      32'H4724: READ <= 8'H61;
      32'H4725: READ <= 8'H5b;
      32'H4726: READ <= 8'H45;
      32'H4727: READ <= 8'H2d;
      32'H4728: READ <= 8'H27;
      32'H4729: READ <= 8'H22;
      32'H4730: READ <= 8'H1d;
      32'H4731: READ <= 8'H1a;
      32'H4732: READ <= 8'H16;
      32'H4733: READ <= 8'He;
      32'H4734: READ <= 8'Ha;
      32'H4735: READ <= 8'H6;
      32'H4736: READ <= 8'H20;
      32'H4737: READ <= 8'H44;
      32'H4738: READ <= 8'H26;
      32'H4739: READ <= 8'H50;
      32'H4740: READ <= 8'H1e;
      32'H4741: READ <= 8'H15;
      32'H4742: READ <= 8'H26;
      32'H4743: READ <= 8'H3a;
      32'H4744: READ <= 8'Hbb;
      32'H4745: READ <= 8'Hea;
      32'H4746: READ <= 8'Hea;
      32'H4747: READ <= 8'He5;
      32'H4748: READ <= 8'He6;
      32'H4749: READ <= 8'He0;
      32'H4750: READ <= 8'Hd2;
      32'H4751: READ <= 8'Hc5;
      32'H4752: READ <= 8'Hb9;
      32'H4753: READ <= 8'Ha5;
      32'H4754: READ <= 8'Ha8;
      32'H4755: READ <= 8'Ha4;
      32'H4756: READ <= 8'H8e;
      32'H4757: READ <= 8'H7a;
      32'H4758: READ <= 8'H74;
      32'H4759: READ <= 8'H3a;
      32'H4760: READ <= 8'H34;
      32'H4761: READ <= 8'H7c;
      32'H4762: READ <= 8'H74;
      32'H4763: READ <= 8'H72;
      32'H4764: READ <= 8'H3a;
      32'H4765: READ <= 8'H5d;
      32'H4766: READ <= 8'H62;
      32'H4767: READ <= 8'H64;
      32'H4768: READ <= 8'H73;
      32'H4769: READ <= 8'H77;
      32'H4770: READ <= 8'H81;
      32'H4771: READ <= 8'H83;
      32'H4772: READ <= 8'H84;
      32'H4773: READ <= 8'H90;
      32'H4774: READ <= 8'H9a;
      32'H4775: READ <= 8'H9e;
      32'H4776: READ <= 8'Hb1;
      32'H4777: READ <= 8'H98;
      32'H4778: READ <= 8'H88;
      32'H4779: READ <= 8'H7b;
      32'H4780: READ <= 8'H7b;
      32'H4781: READ <= 8'H7b;
      32'H4782: READ <= 8'H7c;
      32'H4783: READ <= 8'H7d;
      32'H4784: READ <= 8'H7d;
      32'H4785: READ <= 8'H7f;
      32'H4786: READ <= 8'H81;
      32'H4787: READ <= 8'H81;
      32'H4788: READ <= 8'H82;
      32'H4789: READ <= 8'H83;
      32'H4790: READ <= 8'H84;
      32'H4791: READ <= 8'H85;
      32'H4792: READ <= 8'H86;
      32'H4793: READ <= 8'H87;
      32'H4794: READ <= 8'H88;
      32'H4795: READ <= 8'H88;
      32'H4796: READ <= 8'H89;
      32'H4797: READ <= 8'H89;
      32'H4798: READ <= 8'H89;
      32'H4799: READ <= 8'H8a;
      32'H4800: READ <= 8'H71;
      32'H4801: READ <= 8'H71;
      32'H4802: READ <= 8'H71;
      32'H4803: READ <= 8'H70;
      32'H4804: READ <= 8'H71;
      32'H4805: READ <= 8'H71;
      32'H4806: READ <= 8'H72;
      32'H4807: READ <= 8'H73;
      32'H4808: READ <= 8'H73;
      32'H4809: READ <= 8'H72;
      32'H4810: READ <= 8'H72;
      32'H4811: READ <= 8'H72;
      32'H4812: READ <= 8'H72;
      32'H4813: READ <= 8'H73;
      32'H4814: READ <= 8'H73;
      32'H4815: READ <= 8'H74;
      32'H4816: READ <= 8'H75;
      32'H4817: READ <= 8'H77;
      32'H4818: READ <= 8'H82;
      32'H4819: READ <= 8'H90;
      32'H4820: READ <= 8'Had;
      32'H4821: READ <= 8'Hbe;
      32'H4822: READ <= 8'Hbc;
      32'H4823: READ <= 8'H99;
      32'H4824: READ <= 8'H65;
      32'H4825: READ <= 8'H60;
      32'H4826: READ <= 8'H51;
      32'H4827: READ <= 8'H22;
      32'H4828: READ <= 8'H20;
      32'H4829: READ <= 8'H1f;
      32'H4830: READ <= 8'H1e;
      32'H4831: READ <= 8'H1c;
      32'H4832: READ <= 8'H18;
      32'H4833: READ <= 8'Hf;
      32'H4834: READ <= 8'H9;
      32'H4835: READ <= 8'H7;
      32'H4836: READ <= 8'He;
      32'H4837: READ <= 8'H48;
      32'H4838: READ <= 8'H2e;
      32'H4839: READ <= 8'H4c;
      32'H4840: READ <= 8'H44;
      32'H4841: READ <= 8'H21;
      32'H4842: READ <= 8'H33;
      32'H4843: READ <= 8'H8f;
      32'H4844: READ <= 8'He1;
      32'H4845: READ <= 8'He2;
      32'H4846: READ <= 8'Hdb;
      32'H4847: READ <= 8'Hd8;
      32'H4848: READ <= 8'Hdf;
      32'H4849: READ <= 8'He2;
      32'H4850: READ <= 8'Hdd;
      32'H4851: READ <= 8'Hdc;
      32'H4852: READ <= 8'Hcc;
      32'H4853: READ <= 8'Hb0;
      32'H4854: READ <= 8'Ha1;
      32'H4855: READ <= 8'Ha3;
      32'H4856: READ <= 8'H9e;
      32'H4857: READ <= 8'H86;
      32'H4858: READ <= 8'H8e;
      32'H4859: READ <= 8'H37;
      32'H4860: READ <= 8'H5a;
      32'H4861: READ <= 8'H87;
      32'H4862: READ <= 8'H8c;
      32'H4863: READ <= 8'H71;
      32'H4864: READ <= 8'H34;
      32'H4865: READ <= 8'H62;
      32'H4866: READ <= 8'H64;
      32'H4867: READ <= 8'H71;
      32'H4868: READ <= 8'H66;
      32'H4869: READ <= 8'H75;
      32'H4870: READ <= 8'H80;
      32'H4871: READ <= 8'H81;
      32'H4872: READ <= 8'H85;
      32'H4873: READ <= 8'H99;
      32'H4874: READ <= 8'H9d;
      32'H4875: READ <= 8'Hab;
      32'H4876: READ <= 8'Haa;
      32'H4877: READ <= 8'H90;
      32'H4878: READ <= 8'H81;
      32'H4879: READ <= 8'H7b;
      32'H4880: READ <= 8'H7b;
      32'H4881: READ <= 8'H7b;
      32'H4882: READ <= 8'H7c;
      32'H4883: READ <= 8'H7d;
      32'H4884: READ <= 8'H7e;
      32'H4885: READ <= 8'H7f;
      32'H4886: READ <= 8'H80;
      32'H4887: READ <= 8'H81;
      32'H4888: READ <= 8'H82;
      32'H4889: READ <= 8'H83;
      32'H4890: READ <= 8'H84;
      32'H4891: READ <= 8'H85;
      32'H4892: READ <= 8'H86;
      32'H4893: READ <= 8'H87;
      32'H4894: READ <= 8'H89;
      32'H4895: READ <= 8'H88;
      32'H4896: READ <= 8'H89;
      32'H4897: READ <= 8'H89;
      32'H4898: READ <= 8'H8a;
      32'H4899: READ <= 8'H8a;
      32'H4900: READ <= 8'H70;
      32'H4901: READ <= 8'H70;
      32'H4902: READ <= 8'H70;
      32'H4903: READ <= 8'H70;
      32'H4904: READ <= 8'H70;
      32'H4905: READ <= 8'H71;
      32'H4906: READ <= 8'H71;
      32'H4907: READ <= 8'H71;
      32'H4908: READ <= 8'H72;
      32'H4909: READ <= 8'H72;
      32'H4910: READ <= 8'H72;
      32'H4911: READ <= 8'H71;
      32'H4912: READ <= 8'H71;
      32'H4913: READ <= 8'H71;
      32'H4914: READ <= 8'H72;
      32'H4915: READ <= 8'H73;
      32'H4916: READ <= 8'H74;
      32'H4917: READ <= 8'H76;
      32'H4918: READ <= 8'H79;
      32'H4919: READ <= 8'H7f;
      32'H4920: READ <= 8'H97;
      32'H4921: READ <= 8'Had;
      32'H4922: READ <= 8'Hb7;
      32'H4923: READ <= 8'Hb7;
      32'H4924: READ <= 8'H91;
      32'H4925: READ <= 8'H69;
      32'H4926: READ <= 8'H66;
      32'H4927: READ <= 8'H3c;
      32'H4928: READ <= 8'H1e;
      32'H4929: READ <= 8'H1c;
      32'H4930: READ <= 8'H20;
      32'H4931: READ <= 8'H20;
      32'H4932: READ <= 8'H19;
      32'H4933: READ <= 8'He;
      32'H4934: READ <= 8'H8;
      32'H4935: READ <= 8'H6;
      32'H4936: READ <= 8'Hb;
      32'H4937: READ <= 8'H40;
      32'H4938: READ <= 8'H34;
      32'H4939: READ <= 8'H50;
      32'H4940: READ <= 8'H75;
      32'H4941: READ <= 8'H3c;
      32'H4942: READ <= 8'H51;
      32'H4943: READ <= 8'Hc6;
      32'H4944: READ <= 8'Hcd;
      32'H4945: READ <= 8'Hd6;
      32'H4946: READ <= 8'Hd8;
      32'H4947: READ <= 8'Hdb;
      32'H4948: READ <= 8'Hde;
      32'H4949: READ <= 8'Hdb;
      32'H4950: READ <= 8'Hd8;
      32'H4951: READ <= 8'Hd6;
      32'H4952: READ <= 8'Hc6;
      32'H4953: READ <= 8'Hb3;
      32'H4954: READ <= 8'Ha8;
      32'H4955: READ <= 8'H9e;
      32'H4956: READ <= 8'H9a;
      32'H4957: READ <= 8'H8b;
      32'H4958: READ <= 8'H9a;
      32'H4959: READ <= 8'H45;
      32'H4960: READ <= 8'H65;
      32'H4961: READ <= 8'H9b;
      32'H4962: READ <= 8'H89;
      32'H4963: READ <= 8'H8c;
      32'H4964: READ <= 8'H35;
      32'H4965: READ <= 8'H4f;
      32'H4966: READ <= 8'H59;
      32'H4967: READ <= 8'H60;
      32'H4968: READ <= 8'H63;
      32'H4969: READ <= 8'H6f;
      32'H4970: READ <= 8'H73;
      32'H4971: READ <= 8'H83;
      32'H4972: READ <= 8'H89;
      32'H4973: READ <= 8'H99;
      32'H4974: READ <= 8'H9d;
      32'H4975: READ <= 8'Ha2;
      32'H4976: READ <= 8'H8e;
      32'H4977: READ <= 8'H84;
      32'H4978: READ <= 8'H7a;
      32'H4979: READ <= 8'H7b;
      32'H4980: READ <= 8'H7b;
      32'H4981: READ <= 8'H7c;
      32'H4982: READ <= 8'H7d;
      32'H4983: READ <= 8'H7d;
      32'H4984: READ <= 8'H7e;
      32'H4985: READ <= 8'H7f;
      32'H4986: READ <= 8'H80;
      32'H4987: READ <= 8'H81;
      32'H4988: READ <= 8'H82;
      32'H4989: READ <= 8'H82;
      32'H4990: READ <= 8'H84;
      32'H4991: READ <= 8'H84;
      32'H4992: READ <= 8'H86;
      32'H4993: READ <= 8'H87;
      32'H4994: READ <= 8'H88;
      32'H4995: READ <= 8'H88;
      32'H4996: READ <= 8'H89;
      32'H4997: READ <= 8'H89;
      32'H4998: READ <= 8'H8a;
      32'H4999: READ <= 8'H8a;
      32'H5000: READ <= 8'H70;
      32'H5001: READ <= 8'H70;
      32'H5002: READ <= 8'H70;
      32'H5003: READ <= 8'H70;
      32'H5004: READ <= 8'H6f;
      32'H5005: READ <= 8'H70;
      32'H5006: READ <= 8'H70;
      32'H5007: READ <= 8'H70;
      32'H5008: READ <= 8'H71;
      32'H5009: READ <= 8'H71;
      32'H5010: READ <= 8'H71;
      32'H5011: READ <= 8'H71;
      32'H5012: READ <= 8'H70;
      32'H5013: READ <= 8'H71;
      32'H5014: READ <= 8'H71;
      32'H5015: READ <= 8'H72;
      32'H5016: READ <= 8'H73;
      32'H5017: READ <= 8'H74;
      32'H5018: READ <= 8'H77;
      32'H5019: READ <= 8'H78;
      32'H5020: READ <= 8'H87;
      32'H5021: READ <= 8'H8e;
      32'H5022: READ <= 8'H97;
      32'H5023: READ <= 8'H96;
      32'H5024: READ <= 8'Ha0;
      32'H5025: READ <= 8'H8f;
      32'H5026: READ <= 8'H84;
      32'H5027: READ <= 8'H77;
      32'H5028: READ <= 8'H4a;
      32'H5029: READ <= 8'H2f;
      32'H5030: READ <= 8'H2a;
      32'H5031: READ <= 8'H27;
      32'H5032: READ <= 8'H1d;
      32'H5033: READ <= 8'H13;
      32'H5034: READ <= 8'Hf;
      32'H5035: READ <= 8'Hc;
      32'H5036: READ <= 8'Hc;
      32'H5037: READ <= 8'H2c;
      32'H5038: READ <= 8'H29;
      32'H5039: READ <= 8'H54;
      32'H5040: READ <= 8'H4d;
      32'H5041: READ <= 8'H61;
      32'H5042: READ <= 8'H85;
      32'H5043: READ <= 8'Hb2;
      32'H5044: READ <= 8'Hb9;
      32'H5045: READ <= 8'Hd4;
      32'H5046: READ <= 8'Hde;
      32'H5047: READ <= 8'He2;
      32'H5048: READ <= 8'He7;
      32'H5049: READ <= 8'He6;
      32'H5050: READ <= 8'He0;
      32'H5051: READ <= 8'Hd9;
      32'H5052: READ <= 8'Hc9;
      32'H5053: READ <= 8'Had;
      32'H5054: READ <= 8'Hb2;
      32'H5055: READ <= 8'H9b;
      32'H5056: READ <= 8'H9e;
      32'H5057: READ <= 8'H8f;
      32'H5058: READ <= 8'H9f;
      32'H5059: READ <= 8'H4f;
      32'H5060: READ <= 8'H52;
      32'H5061: READ <= 8'H9f;
      32'H5062: READ <= 8'H78;
      32'H5063: READ <= 8'Ha1;
      32'H5064: READ <= 8'H37;
      32'H5065: READ <= 8'H59;
      32'H5066: READ <= 8'H5d;
      32'H5067: READ <= 8'H6a;
      32'H5068: READ <= 8'H65;
      32'H5069: READ <= 8'H5d;
      32'H5070: READ <= 8'H62;
      32'H5071: READ <= 8'H67;
      32'H5072: READ <= 8'H72;
      32'H5073: READ <= 8'H84;
      32'H5074: READ <= 8'H8e;
      32'H5075: READ <= 8'H91;
      32'H5076: READ <= 8'H92;
      32'H5077: READ <= 8'H7c;
      32'H5078: READ <= 8'H7a;
      32'H5079: READ <= 8'H7a;
      32'H5080: READ <= 8'H7a;
      32'H5081: READ <= 8'H7b;
      32'H5082: READ <= 8'H7c;
      32'H5083: READ <= 8'H7e;
      32'H5084: READ <= 8'H7e;
      32'H5085: READ <= 8'H7f;
      32'H5086: READ <= 8'H80;
      32'H5087: READ <= 8'H81;
      32'H5088: READ <= 8'H82;
      32'H5089: READ <= 8'H83;
      32'H5090: READ <= 8'H83;
      32'H5091: READ <= 8'H85;
      32'H5092: READ <= 8'H86;
      32'H5093: READ <= 8'H87;
      32'H5094: READ <= 8'H88;
      32'H5095: READ <= 8'H89;
      32'H5096: READ <= 8'H89;
      32'H5097: READ <= 8'H8a;
      32'H5098: READ <= 8'H8a;
      32'H5099: READ <= 8'H89;
      32'H5100: READ <= 8'H70;
      32'H5101: READ <= 8'H6f;
      32'H5102: READ <= 8'H6f;
      32'H5103: READ <= 8'H6f;
      32'H5104: READ <= 8'H70;
      32'H5105: READ <= 8'H70;
      32'H5106: READ <= 8'H70;
      32'H5107: READ <= 8'H6f;
      32'H5108: READ <= 8'H70;
      32'H5109: READ <= 8'H70;
      32'H5110: READ <= 8'H70;
      32'H5111: READ <= 8'H71;
      32'H5112: READ <= 8'H6f;
      32'H5113: READ <= 8'H6f;
      32'H5114: READ <= 8'H70;
      32'H5115: READ <= 8'H71;
      32'H5116: READ <= 8'H72;
      32'H5117: READ <= 8'H74;
      32'H5118: READ <= 8'H76;
      32'H5119: READ <= 8'H78;
      32'H5120: READ <= 8'H7b;
      32'H5121: READ <= 8'H7d;
      32'H5122: READ <= 8'H82;
      32'H5123: READ <= 8'H87;
      32'H5124: READ <= 8'H8c;
      32'H5125: READ <= 8'H92;
      32'H5126: READ <= 8'H9e;
      32'H5127: READ <= 8'H8c;
      32'H5128: READ <= 8'H5d;
      32'H5129: READ <= 8'H4f;
      32'H5130: READ <= 8'H45;
      32'H5131: READ <= 8'H40;
      32'H5132: READ <= 8'H31;
      32'H5133: READ <= 8'H24;
      32'H5134: READ <= 8'H19;
      32'H5135: READ <= 8'Hf;
      32'H5136: READ <= 8'H1f;
      32'H5137: READ <= 8'H37;
      32'H5138: READ <= 8'H34;
      32'H5139: READ <= 8'H28;
      32'H5140: READ <= 8'H29;
      32'H5141: READ <= 8'H70;
      32'H5142: READ <= 8'H8d;
      32'H5143: READ <= 8'Ha2;
      32'H5144: READ <= 8'Hc1;
      32'H5145: READ <= 8'Hda;
      32'H5146: READ <= 8'He0;
      32'H5147: READ <= 8'He4;
      32'H5148: READ <= 8'He9;
      32'H5149: READ <= 8'Heb;
      32'H5150: READ <= 8'He8;
      32'H5151: READ <= 8'He1;
      32'H5152: READ <= 8'Hd1;
      32'H5153: READ <= 8'Hbc;
      32'H5154: READ <= 8'Hbe;
      32'H5155: READ <= 8'Hb2;
      32'H5156: READ <= 8'H9a;
      32'H5157: READ <= 8'H9d;
      32'H5158: READ <= 8'H9b;
      32'H5159: READ <= 8'H61;
      32'H5160: READ <= 8'H47;
      32'H5161: READ <= 8'Ha1;
      32'H5162: READ <= 8'H75;
      32'H5163: READ <= 8'H9b;
      32'H5164: READ <= 8'H4a;
      32'H5165: READ <= 8'H7a;
      32'H5166: READ <= 8'H64;
      32'H5167: READ <= 8'H64;
      32'H5168: READ <= 8'H70;
      32'H5169: READ <= 8'H73;
      32'H5170: READ <= 8'H7f;
      32'H5171: READ <= 8'H85;
      32'H5172: READ <= 8'H91;
      32'H5173: READ <= 8'Ha0;
      32'H5174: READ <= 8'Ha8;
      32'H5175: READ <= 8'Ha1;
      32'H5176: READ <= 8'H91;
      32'H5177: READ <= 8'H78;
      32'H5178: READ <= 8'H7a;
      32'H5179: READ <= 8'H7a;
      32'H5180: READ <= 8'H7a;
      32'H5181: READ <= 8'H7b;
      32'H5182: READ <= 8'H7d;
      32'H5183: READ <= 8'H7e;
      32'H5184: READ <= 8'H7e;
      32'H5185: READ <= 8'H7f;
      32'H5186: READ <= 8'H80;
      32'H5187: READ <= 8'H81;
      32'H5188: READ <= 8'H81;
      32'H5189: READ <= 8'H83;
      32'H5190: READ <= 8'H83;
      32'H5191: READ <= 8'H84;
      32'H5192: READ <= 8'H86;
      32'H5193: READ <= 8'H87;
      32'H5194: READ <= 8'H88;
      32'H5195: READ <= 8'H89;
      32'H5196: READ <= 8'H89;
      32'H5197: READ <= 8'H8a;
      32'H5198: READ <= 8'H8a;
      32'H5199: READ <= 8'H89;
      32'H5200: READ <= 8'H70;
      32'H5201: READ <= 8'H70;
      32'H5202: READ <= 8'H6f;
      32'H5203: READ <= 8'H6f;
      32'H5204: READ <= 8'H6f;
      32'H5205: READ <= 8'H6f;
      32'H5206: READ <= 8'H6f;
      32'H5207: READ <= 8'H6f;
      32'H5208: READ <= 8'H6f;
      32'H5209: READ <= 8'H70;
      32'H5210: READ <= 8'H6f;
      32'H5211: READ <= 8'H6f;
      32'H5212: READ <= 8'H6f;
      32'H5213: READ <= 8'H6f;
      32'H5214: READ <= 8'H6f;
      32'H5215: READ <= 8'H70;
      32'H5216: READ <= 8'H71;
      32'H5217: READ <= 8'H72;
      32'H5218: READ <= 8'H73;
      32'H5219: READ <= 8'H77;
      32'H5220: READ <= 8'H78;
      32'H5221: READ <= 8'H7a;
      32'H5222: READ <= 8'H7e;
      32'H5223: READ <= 8'H81;
      32'H5224: READ <= 8'H86;
      32'H5225: READ <= 8'H91;
      32'H5226: READ <= 8'H8b;
      32'H5227: READ <= 8'H57;
      32'H5228: READ <= 8'H55;
      32'H5229: READ <= 8'H57;
      32'H5230: READ <= 8'H31;
      32'H5231: READ <= 8'H1a;
      32'H5232: READ <= 8'H1f;
      32'H5233: READ <= 8'H12;
      32'H5234: READ <= 8'Hf;
      32'H5235: READ <= 8'H12;
      32'H5236: READ <= 8'H16;
      32'H5237: READ <= 8'H3f;
      32'H5238: READ <= 8'H2d;
      32'H5239: READ <= 8'H10;
      32'H5240: READ <= 8'H56;
      32'H5241: READ <= 8'H72;
      32'H5242: READ <= 8'H9c;
      32'H5243: READ <= 8'Hb7;
      32'H5244: READ <= 8'Hce;
      32'H5245: READ <= 8'Hde;
      32'H5246: READ <= 8'He2;
      32'H5247: READ <= 8'He5;
      32'H5248: READ <= 8'He9;
      32'H5249: READ <= 8'Heb;
      32'H5250: READ <= 8'He9;
      32'H5251: READ <= 8'He3;
      32'H5252: READ <= 8'Hd1;
      32'H5253: READ <= 8'Hc4;
      32'H5254: READ <= 8'Hc9;
      32'H5255: READ <= 8'Hb7;
      32'H5256: READ <= 8'Ha6;
      32'H5257: READ <= 8'H8c;
      32'H5258: READ <= 8'H90;
      32'H5259: READ <= 8'H71;
      32'H5260: READ <= 8'H33;
      32'H5261: READ <= 8'H9a;
      32'H5262: READ <= 8'H7c;
      32'H5263: READ <= 8'H98;
      32'H5264: READ <= 8'H52;
      32'H5265: READ <= 8'H78;
      32'H5266: READ <= 8'H6c;
      32'H5267: READ <= 8'H65;
      32'H5268: READ <= 8'H77;
      32'H5269: READ <= 8'H87;
      32'H5270: READ <= 8'H83;
      32'H5271: READ <= 8'H9a;
      32'H5272: READ <= 8'Ha2;
      32'H5273: READ <= 8'Ha8;
      32'H5274: READ <= 8'Hb1;
      32'H5275: READ <= 8'Ha5;
      32'H5276: READ <= 8'H7c;
      32'H5277: READ <= 8'H79;
      32'H5278: READ <= 8'H79;
      32'H5279: READ <= 8'H7a;
      32'H5280: READ <= 8'H7b;
      32'H5281: READ <= 8'H7b;
      32'H5282: READ <= 8'H7c;
      32'H5283: READ <= 8'H7d;
      32'H5284: READ <= 8'H7e;
      32'H5285: READ <= 8'H7f;
      32'H5286: READ <= 8'H80;
      32'H5287: READ <= 8'H80;
      32'H5288: READ <= 8'H81;
      32'H5289: READ <= 8'H82;
      32'H5290: READ <= 8'H84;
      32'H5291: READ <= 8'H85;
      32'H5292: READ <= 8'H86;
      32'H5293: READ <= 8'H87;
      32'H5294: READ <= 8'H87;
      32'H5295: READ <= 8'H89;
      32'H5296: READ <= 8'H89;
      32'H5297: READ <= 8'H89;
      32'H5298: READ <= 8'H8a;
      32'H5299: READ <= 8'H8a;
      32'H5300: READ <= 8'H70;
      32'H5301: READ <= 8'H70;
      32'H5302: READ <= 8'H6f;
      32'H5303: READ <= 8'H70;
      32'H5304: READ <= 8'H6f;
      32'H5305: READ <= 8'H6f;
      32'H5306: READ <= 8'H6e;
      32'H5307: READ <= 8'H6f;
      32'H5308: READ <= 8'H6e;
      32'H5309: READ <= 8'H6e;
      32'H5310: READ <= 8'H6e;
      32'H5311: READ <= 8'H6e;
      32'H5312: READ <= 8'H6e;
      32'H5313: READ <= 8'H6e;
      32'H5314: READ <= 8'H6e;
      32'H5315: READ <= 8'H6f;
      32'H5316: READ <= 8'H70;
      32'H5317: READ <= 8'H71;
      32'H5318: READ <= 8'H73;
      32'H5319: READ <= 8'H74;
      32'H5320: READ <= 8'H76;
      32'H5321: READ <= 8'H78;
      32'H5322: READ <= 8'H7b;
      32'H5323: READ <= 8'H7d;
      32'H5324: READ <= 8'H7f;
      32'H5325: READ <= 8'H85;
      32'H5326: READ <= 8'H65;
      32'H5327: READ <= 8'H45;
      32'H5328: READ <= 8'H52;
      32'H5329: READ <= 8'H32;
      32'H5330: READ <= 8'H5;
      32'H5331: READ <= 8'H9;
      32'H5332: READ <= 8'Hf;
      32'H5333: READ <= 8'Hf;
      32'H5334: READ <= 8'He;
      32'H5335: READ <= 8'Hd;
      32'H5336: READ <= 8'H1f;
      32'H5337: READ <= 8'H47;
      32'H5338: READ <= 8'H3c;
      32'H5339: READ <= 8'H58;
      32'H5340: READ <= 8'H77;
      32'H5341: READ <= 8'H7f;
      32'H5342: READ <= 8'Hb0;
      32'H5343: READ <= 8'Hc7;
      32'H5344: READ <= 8'Hd9;
      32'H5345: READ <= 8'He0;
      32'H5346: READ <= 8'He3;
      32'H5347: READ <= 8'He6;
      32'H5348: READ <= 8'He9;
      32'H5349: READ <= 8'Heb;
      32'H5350: READ <= 8'He9;
      32'H5351: READ <= 8'He2;
      32'H5352: READ <= 8'Hd3;
      32'H5353: READ <= 8'Hc9;
      32'H5354: READ <= 8'Hca;
      32'H5355: READ <= 8'Hb7;
      32'H5356: READ <= 8'Ha7;
      32'H5357: READ <= 8'H91;
      32'H5358: READ <= 8'H85;
      32'H5359: READ <= 8'H73;
      32'H5360: READ <= 8'H2d;
      32'H5361: READ <= 8'H93;
      32'H5362: READ <= 8'H7d;
      32'H5363: READ <= 8'H85;
      32'H5364: READ <= 8'H57;
      32'H5365: READ <= 8'H79;
      32'H5366: READ <= 8'H77;
      32'H5367: READ <= 8'H52;
      32'H5368: READ <= 8'H65;
      32'H5369: READ <= 8'H77;
      32'H5370: READ <= 8'H93;
      32'H5371: READ <= 8'H97;
      32'H5372: READ <= 8'Ha0;
      32'H5373: READ <= 8'Hb3;
      32'H5374: READ <= 8'Haa;
      32'H5375: READ <= 8'H96;
      32'H5376: READ <= 8'H78;
      32'H5377: READ <= 8'H79;
      32'H5378: READ <= 8'H79;
      32'H5379: READ <= 8'H7a;
      32'H5380: READ <= 8'H7b;
      32'H5381: READ <= 8'H7b;
      32'H5382: READ <= 8'H7d;
      32'H5383: READ <= 8'H7d;
      32'H5384: READ <= 8'H7d;
      32'H5385: READ <= 8'H7e;
      32'H5386: READ <= 8'H80;
      32'H5387: READ <= 8'H80;
      32'H5388: READ <= 8'H81;
      32'H5389: READ <= 8'H82;
      32'H5390: READ <= 8'H84;
      32'H5391: READ <= 8'H85;
      32'H5392: READ <= 8'H86;
      32'H5393: READ <= 8'H86;
      32'H5394: READ <= 8'H87;
      32'H5395: READ <= 8'H88;
      32'H5396: READ <= 8'H89;
      32'H5397: READ <= 8'H8a;
      32'H5398: READ <= 8'H8a;
      32'H5399: READ <= 8'H89;
      32'H5400: READ <= 8'H70;
      32'H5401: READ <= 8'H70;
      32'H5402: READ <= 8'H6f;
      32'H5403: READ <= 8'H6f;
      32'H5404: READ <= 8'H6f;
      32'H5405: READ <= 8'H6f;
      32'H5406: READ <= 8'H6e;
      32'H5407: READ <= 8'H6e;
      32'H5408: READ <= 8'H6e;
      32'H5409: READ <= 8'H6e;
      32'H5410: READ <= 8'H6d;
      32'H5411: READ <= 8'H6d;
      32'H5412: READ <= 8'H6d;
      32'H5413: READ <= 8'H6d;
      32'H5414: READ <= 8'H6e;
      32'H5415: READ <= 8'H6e;
      32'H5416: READ <= 8'H6e;
      32'H5417: READ <= 8'H70;
      32'H5418: READ <= 8'H72;
      32'H5419: READ <= 8'H74;
      32'H5420: READ <= 8'H74;
      32'H5421: READ <= 8'H77;
      32'H5422: READ <= 8'H78;
      32'H5423: READ <= 8'H7b;
      32'H5424: READ <= 8'H7c;
      32'H5425: READ <= 8'H81;
      32'H5426: READ <= 8'H5b;
      32'H5427: READ <= 8'H4c;
      32'H5428: READ <= 8'H5e;
      32'H5429: READ <= 8'Hc;
      32'H5430: READ <= 8'Hd;
      32'H5431: READ <= 8'H14;
      32'H5432: READ <= 8'H16;
      32'H5433: READ <= 8'H13;
      32'H5434: READ <= 8'H1a;
      32'H5435: READ <= 8'H1c;
      32'H5436: READ <= 8'H5f;
      32'H5437: READ <= 8'H45;
      32'H5438: READ <= 8'H4d;
      32'H5439: READ <= 8'H5e;
      32'H5440: READ <= 8'H7e;
      32'H5441: READ <= 8'Ha7;
      32'H5442: READ <= 8'Hc1;
      32'H5443: READ <= 8'Hd0;
      32'H5444: READ <= 8'Hdd;
      32'H5445: READ <= 8'He1;
      32'H5446: READ <= 8'He3;
      32'H5447: READ <= 8'He6;
      32'H5448: READ <= 8'He8;
      32'H5449: READ <= 8'He9;
      32'H5450: READ <= 8'He7;
      32'H5451: READ <= 8'He0;
      32'H5452: READ <= 8'Hd5;
      32'H5453: READ <= 8'Hd0;
      32'H5454: READ <= 8'Hcd;
      32'H5455: READ <= 8'Hc6;
      32'H5456: READ <= 8'Hc3;
      32'H5457: READ <= 8'Hb6;
      32'H5458: READ <= 8'H8b;
      32'H5459: READ <= 8'H75;
      32'H5460: READ <= 8'H16;
      32'H5461: READ <= 8'H94;
      32'H5462: READ <= 8'H82;
      32'H5463: READ <= 8'H76;
      32'H5464: READ <= 8'H65;
      32'H5465: READ <= 8'H7c;
      32'H5466: READ <= 8'H64;
      32'H5467: READ <= 8'H70;
      32'H5468: READ <= 8'H78;
      32'H5469: READ <= 8'H87;
      32'H5470: READ <= 8'H8f;
      32'H5471: READ <= 8'H99;
      32'H5472: READ <= 8'Had;
      32'H5473: READ <= 8'Hb0;
      32'H5474: READ <= 8'Ha9;
      32'H5475: READ <= 8'H83;
      32'H5476: READ <= 8'H78;
      32'H5477: READ <= 8'H79;
      32'H5478: READ <= 8'H79;
      32'H5479: READ <= 8'H7a;
      32'H5480: READ <= 8'H7b;
      32'H5481: READ <= 8'H7b;
      32'H5482: READ <= 8'H7c;
      32'H5483: READ <= 8'H7d;
      32'H5484: READ <= 8'H7e;
      32'H5485: READ <= 8'H7f;
      32'H5486: READ <= 8'H80;
      32'H5487: READ <= 8'H81;
      32'H5488: READ <= 8'H81;
      32'H5489: READ <= 8'H82;
      32'H5490: READ <= 8'H83;
      32'H5491: READ <= 8'H84;
      32'H5492: READ <= 8'H85;
      32'H5493: READ <= 8'H87;
      32'H5494: READ <= 8'H88;
      32'H5495: READ <= 8'H89;
      32'H5496: READ <= 8'H89;
      32'H5497: READ <= 8'H89;
      32'H5498: READ <= 8'H89;
      32'H5499: READ <= 8'H8a;
      32'H5500: READ <= 8'H70;
      32'H5501: READ <= 8'H70;
      32'H5502: READ <= 8'H6f;
      32'H5503: READ <= 8'H70;
      32'H5504: READ <= 8'H70;
      32'H5505: READ <= 8'H6f;
      32'H5506: READ <= 8'H6e;
      32'H5507: READ <= 8'H6d;
      32'H5508: READ <= 8'H6e;
      32'H5509: READ <= 8'H6d;
      32'H5510: READ <= 8'H6d;
      32'H5511: READ <= 8'H6d;
      32'H5512: READ <= 8'H6c;
      32'H5513: READ <= 8'H6c;
      32'H5514: READ <= 8'H6d;
      32'H5515: READ <= 8'H6d;
      32'H5516: READ <= 8'H6d;
      32'H5517: READ <= 8'H6f;
      32'H5518: READ <= 8'H70;
      32'H5519: READ <= 8'H72;
      32'H5520: READ <= 8'H74;
      32'H5521: READ <= 8'H74;
      32'H5522: READ <= 8'H76;
      32'H5523: READ <= 8'H78;
      32'H5524: READ <= 8'H7a;
      32'H5525: READ <= 8'H7b;
      32'H5526: READ <= 8'H82;
      32'H5527: READ <= 8'H8a;
      32'H5528: READ <= 8'H77;
      32'H5529: READ <= 8'H2f;
      32'H5530: READ <= 8'H30;
      32'H5531: READ <= 8'H24;
      32'H5532: READ <= 8'H3f;
      32'H5533: READ <= 8'H62;
      32'H5534: READ <= 8'H7f;
      32'H5535: READ <= 8'H86;
      32'H5536: READ <= 8'H89;
      32'H5537: READ <= 8'H47;
      32'H5538: READ <= 8'H48;
      32'H5539: READ <= 8'H4e;
      32'H5540: READ <= 8'H7e;
      32'H5541: READ <= 8'Hb6;
      32'H5542: READ <= 8'Hc9;
      32'H5543: READ <= 8'Hd5;
      32'H5544: READ <= 8'Hde;
      32'H5545: READ <= 8'He1;
      32'H5546: READ <= 8'He2;
      32'H5547: READ <= 8'He4;
      32'H5548: READ <= 8'He6;
      32'H5549: READ <= 8'He7;
      32'H5550: READ <= 8'He5;
      32'H5551: READ <= 8'Hde;
      32'H5552: READ <= 8'Hd8;
      32'H5553: READ <= 8'Hd4;
      32'H5554: READ <= 8'Hd4;
      32'H5555: READ <= 8'Hd3;
      32'H5556: READ <= 8'Hd3;
      32'H5557: READ <= 8'Hd4;
      32'H5558: READ <= 8'H9e;
      32'H5559: READ <= 8'H71;
      32'H5560: READ <= 8'H17;
      32'H5561: READ <= 8'H7e;
      32'H5562: READ <= 8'H87;
      32'H5563: READ <= 8'H6c;
      32'H5564: READ <= 8'H6e;
      32'H5565: READ <= 8'H73;
      32'H5566: READ <= 8'H6c;
      32'H5567: READ <= 8'H71;
      32'H5568: READ <= 8'H7d;
      32'H5569: READ <= 8'H8a;
      32'H5570: READ <= 8'H98;
      32'H5571: READ <= 8'H9b;
      32'H5572: READ <= 8'Hb1;
      32'H5573: READ <= 8'Haf;
      32'H5574: READ <= 8'H96;
      32'H5575: READ <= 8'H7c;
      32'H5576: READ <= 8'H78;
      32'H5577: READ <= 8'H78;
      32'H5578: READ <= 8'H7a;
      32'H5579: READ <= 8'H7a;
      32'H5580: READ <= 8'H7a;
      32'H5581: READ <= 8'H7b;
      32'H5582: READ <= 8'H7c;
      32'H5583: READ <= 8'H7d;
      32'H5584: READ <= 8'H7e;
      32'H5585: READ <= 8'H7e;
      32'H5586: READ <= 8'H80;
      32'H5587: READ <= 8'H81;
      32'H5588: READ <= 8'H82;
      32'H5589: READ <= 8'H82;
      32'H5590: READ <= 8'H84;
      32'H5591: READ <= 8'H84;
      32'H5592: READ <= 8'H86;
      32'H5593: READ <= 8'H87;
      32'H5594: READ <= 8'H88;
      32'H5595: READ <= 8'H89;
      32'H5596: READ <= 8'H88;
      32'H5597: READ <= 8'H89;
      32'H5598: READ <= 8'H8a;
      32'H5599: READ <= 8'H8a;
      32'H5600: READ <= 8'H70;
      32'H5601: READ <= 8'H70;
      32'H5602: READ <= 8'H70;
      32'H5603: READ <= 8'H6f;
      32'H5604: READ <= 8'H6f;
      32'H5605: READ <= 8'H6e;
      32'H5606: READ <= 8'H6e;
      32'H5607: READ <= 8'H6d;
      32'H5608: READ <= 8'H6d;
      32'H5609: READ <= 8'H6d;
      32'H5610: READ <= 8'H6d;
      32'H5611: READ <= 8'H6c;
      32'H5612: READ <= 8'H6c;
      32'H5613: READ <= 8'H6c;
      32'H5614: READ <= 8'H6c;
      32'H5615: READ <= 8'H6c;
      32'H5616: READ <= 8'H6c;
      32'H5617: READ <= 8'H6d;
      32'H5618: READ <= 8'H6e;
      32'H5619: READ <= 8'H6f;
      32'H5620: READ <= 8'H72;
      32'H5621: READ <= 8'H73;
      32'H5622: READ <= 8'H74;
      32'H5623: READ <= 8'H76;
      32'H5624: READ <= 8'H78;
      32'H5625: READ <= 8'H79;
      32'H5626: READ <= 8'H7c;
      32'H5627: READ <= 8'H7f;
      32'H5628: READ <= 8'H86;
      32'H5629: READ <= 8'H5b;
      32'H5630: READ <= 8'H64;
      32'H5631: READ <= 8'H79;
      32'H5632: READ <= 8'H96;
      32'H5633: READ <= 8'H8e;
      32'H5634: READ <= 8'H8f;
      32'H5635: READ <= 8'H74;
      32'H5636: READ <= 8'H84;
      32'H5637: READ <= 8'H46;
      32'H5638: READ <= 8'H52;
      32'H5639: READ <= 8'H52;
      32'H5640: READ <= 8'H83;
      32'H5641: READ <= 8'Hb7;
      32'H5642: READ <= 8'Hca;
      32'H5643: READ <= 8'Hd5;
      32'H5644: READ <= 8'Hdc;
      32'H5645: READ <= 8'Hdd;
      32'H5646: READ <= 8'Hde;
      32'H5647: READ <= 8'Hdf;
      32'H5648: READ <= 8'He2;
      32'H5649: READ <= 8'He2;
      32'H5650: READ <= 8'He0;
      32'H5651: READ <= 8'Hdd;
      32'H5652: READ <= 8'Hda;
      32'H5653: READ <= 8'Hd9;
      32'H5654: READ <= 8'Hdc;
      32'H5655: READ <= 8'Hde;
      32'H5656: READ <= 8'He3;
      32'H5657: READ <= 8'He3;
      32'H5658: READ <= 8'Hc1;
      32'H5659: READ <= 8'H6e;
      32'H5660: READ <= 8'H18;
      32'H5661: READ <= 8'H79;
      32'H5662: READ <= 8'H85;
      32'H5663: READ <= 8'H6f;
      32'H5664: READ <= 8'H63;
      32'H5665: READ <= 8'H77;
      32'H5666: READ <= 8'H71;
      32'H5667: READ <= 8'H75;
      32'H5668: READ <= 8'H80;
      32'H5669: READ <= 8'H91;
      32'H5670: READ <= 8'H9b;
      32'H5671: READ <= 8'Ha7;
      32'H5672: READ <= 8'Haf;
      32'H5673: READ <= 8'Ha3;
      32'H5674: READ <= 8'H8a;
      32'H5675: READ <= 8'H76;
      32'H5676: READ <= 8'H78;
      32'H5677: READ <= 8'H79;
      32'H5678: READ <= 8'H79;
      32'H5679: READ <= 8'H7a;
      32'H5680: READ <= 8'H7a;
      32'H5681: READ <= 8'H7b;
      32'H5682: READ <= 8'H7c;
      32'H5683: READ <= 8'H7d;
      32'H5684: READ <= 8'H7e;
      32'H5685: READ <= 8'H7e;
      32'H5686: READ <= 8'H80;
      32'H5687: READ <= 8'H80;
      32'H5688: READ <= 8'H81;
      32'H5689: READ <= 8'H82;
      32'H5690: READ <= 8'H83;
      32'H5691: READ <= 8'H84;
      32'H5692: READ <= 8'H86;
      32'H5693: READ <= 8'H87;
      32'H5694: READ <= 8'H88;
      32'H5695: READ <= 8'H88;
      32'H5696: READ <= 8'H88;
      32'H5697: READ <= 8'H89;
      32'H5698: READ <= 8'H89;
      32'H5699: READ <= 8'H89;
      32'H5700: READ <= 8'H70;
      32'H5701: READ <= 8'H70;
      32'H5702: READ <= 8'H70;
      32'H5703: READ <= 8'H6f;
      32'H5704: READ <= 8'H6f;
      32'H5705: READ <= 8'H6e;
      32'H5706: READ <= 8'H6e;
      32'H5707: READ <= 8'H6d;
      32'H5708: READ <= 8'H6d;
      32'H5709: READ <= 8'H6d;
      32'H5710: READ <= 8'H6c;
      32'H5711: READ <= 8'H6c;
      32'H5712: READ <= 8'H6b;
      32'H5713: READ <= 8'H6b;
      32'H5714: READ <= 8'H6b;
      32'H5715: READ <= 8'H6b;
      32'H5716: READ <= 8'H6b;
      32'H5717: READ <= 8'H6c;
      32'H5718: READ <= 8'H6d;
      32'H5719: READ <= 8'H6d;
      32'H5720: READ <= 8'H6f;
      32'H5721: READ <= 8'H71;
      32'H5722: READ <= 8'H72;
      32'H5723: READ <= 8'H73;
      32'H5724: READ <= 8'H76;
      32'H5725: READ <= 8'H77;
      32'H5726: READ <= 8'H7a;
      32'H5727: READ <= 8'H7e;
      32'H5728: READ <= 8'H80;
      32'H5729: READ <= 8'H87;
      32'H5730: READ <= 8'H8a;
      32'H5731: READ <= 8'H89;
      32'H5732: READ <= 8'H87;
      32'H5733: READ <= 8'H88;
      32'H5734: READ <= 8'H8c;
      32'H5735: READ <= 8'H96;
      32'H5736: READ <= 8'H75;
      32'H5737: READ <= 8'H5b;
      32'H5738: READ <= 8'H6e;
      32'H5739: READ <= 8'H65;
      32'H5740: READ <= 8'H8f;
      32'H5741: READ <= 8'Hbe;
      32'H5742: READ <= 8'Hcb;
      32'H5743: READ <= 8'Hd3;
      32'H5744: READ <= 8'Hd8;
      32'H5745: READ <= 8'Hd9;
      32'H5746: READ <= 8'Hd9;
      32'H5747: READ <= 8'Hda;
      32'H5748: READ <= 8'Hdd;
      32'H5749: READ <= 8'Hdd;
      32'H5750: READ <= 8'Hdc;
      32'H5751: READ <= 8'Hdc;
      32'H5752: READ <= 8'Hdd;
      32'H5753: READ <= 8'Hdf;
      32'H5754: READ <= 8'He4;
      32'H5755: READ <= 8'He5;
      32'H5756: READ <= 8'He4;
      32'H5757: READ <= 8'Hea;
      32'H5758: READ <= 8'He9;
      32'H5759: READ <= 8'H73;
      32'H5760: READ <= 8'H1b;
      32'H5761: READ <= 8'H73;
      32'H5762: READ <= 8'H8c;
      32'H5763: READ <= 8'H5f;
      32'H5764: READ <= 8'H58;
      32'H5765: READ <= 8'H74;
      32'H5766: READ <= 8'H6e;
      32'H5767: READ <= 8'H7f;
      32'H5768: READ <= 8'H8d;
      32'H5769: READ <= 8'H90;
      32'H5770: READ <= 8'Ha5;
      32'H5771: READ <= 8'Haf;
      32'H5772: READ <= 8'Ha3;
      32'H5773: READ <= 8'H96;
      32'H5774: READ <= 8'H79;
      32'H5775: READ <= 8'H77;
      32'H5776: READ <= 8'H78;
      32'H5777: READ <= 8'H78;
      32'H5778: READ <= 8'H79;
      32'H5779: READ <= 8'H7a;
      32'H5780: READ <= 8'H7a;
      32'H5781: READ <= 8'H7b;
      32'H5782: READ <= 8'H7c;
      32'H5783: READ <= 8'H7d;
      32'H5784: READ <= 8'H7d;
      32'H5785: READ <= 8'H7e;
      32'H5786: READ <= 8'H7f;
      32'H5787: READ <= 8'H80;
      32'H5788: READ <= 8'H80;
      32'H5789: READ <= 8'H82;
      32'H5790: READ <= 8'H83;
      32'H5791: READ <= 8'H85;
      32'H5792: READ <= 8'H86;
      32'H5793: READ <= 8'H86;
      32'H5794: READ <= 8'H87;
      32'H5795: READ <= 8'H88;
      32'H5796: READ <= 8'H88;
      32'H5797: READ <= 8'H88;
      32'H5798: READ <= 8'H89;
      32'H5799: READ <= 8'H8a;
      32'H5800: READ <= 8'H71;
      32'H5801: READ <= 8'H71;
      32'H5802: READ <= 8'H70;
      32'H5803: READ <= 8'H70;
      32'H5804: READ <= 8'H6f;
      32'H5805: READ <= 8'H6f;
      32'H5806: READ <= 8'H6e;
      32'H5807: READ <= 8'H6e;
      32'H5808: READ <= 8'H6d;
      32'H5809: READ <= 8'H6d;
      32'H5810: READ <= 8'H6c;
      32'H5811: READ <= 8'H6b;
      32'H5812: READ <= 8'H6b;
      32'H5813: READ <= 8'H6a;
      32'H5814: READ <= 8'H6b;
      32'H5815: READ <= 8'H6a;
      32'H5816: READ <= 8'H6a;
      32'H5817: READ <= 8'H6b;
      32'H5818: READ <= 8'H6b;
      32'H5819: READ <= 8'H6c;
      32'H5820: READ <= 8'H6d;
      32'H5821: READ <= 8'H6f;
      32'H5822: READ <= 8'H71;
      32'H5823: READ <= 8'H72;
      32'H5824: READ <= 8'H73;
      32'H5825: READ <= 8'H75;
      32'H5826: READ <= 8'H78;
      32'H5827: READ <= 8'H7c;
      32'H5828: READ <= 8'H7e;
      32'H5829: READ <= 8'H80;
      32'H5830: READ <= 8'H83;
      32'H5831: READ <= 8'H85;
      32'H5832: READ <= 8'H87;
      32'H5833: READ <= 8'H88;
      32'H5834: READ <= 8'H94;
      32'H5835: READ <= 8'H94;
      32'H5836: READ <= 8'H55;
      32'H5837: READ <= 8'H84;
      32'H5838: READ <= 8'H85;
      32'H5839: READ <= 8'H70;
      32'H5840: READ <= 8'H9c;
      32'H5841: READ <= 8'Hc9;
      32'H5842: READ <= 8'Hce;
      32'H5843: READ <= 8'Hd2;
      32'H5844: READ <= 8'Hd4;
      32'H5845: READ <= 8'Hd4;
      32'H5846: READ <= 8'Hd3;
      32'H5847: READ <= 8'Hd4;
      32'H5848: READ <= 8'Hd6;
      32'H5849: READ <= 8'Hd7;
      32'H5850: READ <= 8'Hd8;
      32'H5851: READ <= 8'Hdb;
      32'H5852: READ <= 8'Hdf;
      32'H5853: READ <= 8'He3;
      32'H5854: READ <= 8'He8;
      32'H5855: READ <= 8'He8;
      32'H5856: READ <= 8'He2;
      32'H5857: READ <= 8'He1;
      32'H5858: READ <= 8'He7;
      32'H5859: READ <= 8'H79;
      32'H5860: READ <= 8'H24;
      32'H5861: READ <= 8'H7f;
      32'H5862: READ <= 8'H8e;
      32'H5863: READ <= 8'H59;
      32'H5864: READ <= 8'H50;
      32'H5865: READ <= 8'H7f;
      32'H5866: READ <= 8'H7a;
      32'H5867: READ <= 8'H7e;
      32'H5868: READ <= 8'H8f;
      32'H5869: READ <= 8'H9a;
      32'H5870: READ <= 8'Ha8;
      32'H5871: READ <= 8'Ha6;
      32'H5872: READ <= 8'H98;
      32'H5873: READ <= 8'H7a;
      32'H5874: READ <= 8'H76;
      32'H5875: READ <= 8'H77;
      32'H5876: READ <= 8'H78;
      32'H5877: READ <= 8'H78;
      32'H5878: READ <= 8'H79;
      32'H5879: READ <= 8'H7a;
      32'H5880: READ <= 8'H7b;
      32'H5881: READ <= 8'H7b;
      32'H5882: READ <= 8'H7c;
      32'H5883: READ <= 8'H7c;
      32'H5884: READ <= 8'H7d;
      32'H5885: READ <= 8'H7e;
      32'H5886: READ <= 8'H7f;
      32'H5887: READ <= 8'H80;
      32'H5888: READ <= 8'H81;
      32'H5889: READ <= 8'H83;
      32'H5890: READ <= 8'H83;
      32'H5891: READ <= 8'H84;
      32'H5892: READ <= 8'H86;
      32'H5893: READ <= 8'H86;
      32'H5894: READ <= 8'H87;
      32'H5895: READ <= 8'H88;
      32'H5896: READ <= 8'H88;
      32'H5897: READ <= 8'H88;
      32'H5898: READ <= 8'H89;
      32'H5899: READ <= 8'H89;
      32'H5900: READ <= 8'H72;
      32'H5901: READ <= 8'H71;
      32'H5902: READ <= 8'H71;
      32'H5903: READ <= 8'H71;
      32'H5904: READ <= 8'H70;
      32'H5905: READ <= 8'H6f;
      32'H5906: READ <= 8'H6e;
      32'H5907: READ <= 8'H6e;
      32'H5908: READ <= 8'H6e;
      32'H5909: READ <= 8'H6d;
      32'H5910: READ <= 8'H6d;
      32'H5911: READ <= 8'H6b;
      32'H5912: READ <= 8'H6b;
      32'H5913: READ <= 8'H6a;
      32'H5914: READ <= 8'H6a;
      32'H5915: READ <= 8'H69;
      32'H5916: READ <= 8'H69;
      32'H5917: READ <= 8'H69;
      32'H5918: READ <= 8'H6a;
      32'H5919: READ <= 8'H6b;
      32'H5920: READ <= 8'H6c;
      32'H5921: READ <= 8'H6c;
      32'H5922: READ <= 8'H6e;
      32'H5923: READ <= 8'H71;
      32'H5924: READ <= 8'H72;
      32'H5925: READ <= 8'H74;
      32'H5926: READ <= 8'H76;
      32'H5927: READ <= 8'H7a;
      32'H5928: READ <= 8'H7d;
      32'H5929: READ <= 8'H80;
      32'H5930: READ <= 8'H83;
      32'H5931: READ <= 8'H87;
      32'H5932: READ <= 8'H8a;
      32'H5933: READ <= 8'H8c;
      32'H5934: READ <= 8'H9c;
      32'H5935: READ <= 8'H7e;
      32'H5936: READ <= 8'H5d;
      32'H5937: READ <= 8'H84;
      32'H5938: READ <= 8'H85;
      32'H5939: READ <= 8'H7a;
      32'H5940: READ <= 8'Hb4;
      32'H5941: READ <= 8'Hd6;
      32'H5942: READ <= 8'Hd2;
      32'H5943: READ <= 8'Hd0;
      32'H5944: READ <= 8'Hd0;
      32'H5945: READ <= 8'Hd0;
      32'H5946: READ <= 8'Hd1;
      32'H5947: READ <= 8'Hd1;
      32'H5948: READ <= 8'Hd2;
      32'H5949: READ <= 8'Hd3;
      32'H5950: READ <= 8'Hd6;
      32'H5951: READ <= 8'Hdb;
      32'H5952: READ <= 8'He0;
      32'H5953: READ <= 8'He5;
      32'H5954: READ <= 8'Hea;
      32'H5955: READ <= 8'Heb;
      32'H5956: READ <= 8'He6;
      32'H5957: READ <= 8'He5;
      32'H5958: READ <= 8'He4;
      32'H5959: READ <= 8'H98;
      32'H5960: READ <= 8'H27;
      32'H5961: READ <= 8'H7c;
      32'H5962: READ <= 8'H7d;
      32'H5963: READ <= 8'H5a;
      32'H5964: READ <= 8'H4c;
      32'H5965: READ <= 8'H89;
      32'H5966: READ <= 8'H72;
      32'H5967: READ <= 8'H90;
      32'H5968: READ <= 8'H95;
      32'H5969: READ <= 8'Ha3;
      32'H5970: READ <= 8'Ha0;
      32'H5971: READ <= 8'H98;
      32'H5972: READ <= 8'H8f;
      32'H5973: READ <= 8'H71;
      32'H5974: READ <= 8'H75;
      32'H5975: READ <= 8'H76;
      32'H5976: READ <= 8'H78;
      32'H5977: READ <= 8'H78;
      32'H5978: READ <= 8'H79;
      32'H5979: READ <= 8'H7a;
      32'H5980: READ <= 8'H7a;
      32'H5981: READ <= 8'H7b;
      32'H5982: READ <= 8'H7c;
      32'H5983: READ <= 8'H7c;
      32'H5984: READ <= 8'H7d;
      32'H5985: READ <= 8'H7e;
      32'H5986: READ <= 8'H7f;
      32'H5987: READ <= 8'H80;
      32'H5988: READ <= 8'H81;
      32'H5989: READ <= 8'H82;
      32'H5990: READ <= 8'H83;
      32'H5991: READ <= 8'H84;
      32'H5992: READ <= 8'H85;
      32'H5993: READ <= 8'H86;
      32'H5994: READ <= 8'H87;
      32'H5995: READ <= 8'H87;
      32'H5996: READ <= 8'H88;
      32'H5997: READ <= 8'H88;
      32'H5998: READ <= 8'H89;
      32'H5999: READ <= 8'H8a;
      32'H6000: READ <= 8'H71;
      32'H6001: READ <= 8'H71;
      32'H6002: READ <= 8'H71;
      32'H6003: READ <= 8'H71;
      32'H6004: READ <= 8'H70;
      32'H6005: READ <= 8'H70;
      32'H6006: READ <= 8'H6f;
      32'H6007: READ <= 8'H6e;
      32'H6008: READ <= 8'H6e;
      32'H6009: READ <= 8'H6d;
      32'H6010: READ <= 8'H6d;
      32'H6011: READ <= 8'H6c;
      32'H6012: READ <= 8'H6c;
      32'H6013: READ <= 8'H6b;
      32'H6014: READ <= 8'H6a;
      32'H6015: READ <= 8'H6a;
      32'H6016: READ <= 8'H69;
      32'H6017: READ <= 8'H69;
      32'H6018: READ <= 8'H68;
      32'H6019: READ <= 8'H68;
      32'H6020: READ <= 8'H6a;
      32'H6021: READ <= 8'H6a;
      32'H6022: READ <= 8'H6c;
      32'H6023: READ <= 8'H6e;
      32'H6024: READ <= 8'H70;
      32'H6025: READ <= 8'H73;
      32'H6026: READ <= 8'H76;
      32'H6027: READ <= 8'H79;
      32'H6028: READ <= 8'H7c;
      32'H6029: READ <= 8'H81;
      32'H6030: READ <= 8'H86;
      32'H6031: READ <= 8'H8a;
      32'H6032: READ <= 8'H8d;
      32'H6033: READ <= 8'H91;
      32'H6034: READ <= 8'H99;
      32'H6035: READ <= 8'H5a;
      32'H6036: READ <= 8'Ha6;
      32'H6037: READ <= 8'H8e;
      32'H6038: READ <= 8'H90;
      32'H6039: READ <= 8'H73;
      32'H6040: READ <= 8'Hca;
      32'H6041: READ <= 8'Hd9;
      32'H6042: READ <= 8'Hd4;
      32'H6043: READ <= 8'Hd1;
      32'H6044: READ <= 8'Hce;
      32'H6045: READ <= 8'Hce;
      32'H6046: READ <= 8'Hd1;
      32'H6047: READ <= 8'Hd0;
      32'H6048: READ <= 8'Hd0;
      32'H6049: READ <= 8'Hd1;
      32'H6050: READ <= 8'Hd5;
      32'H6051: READ <= 8'Hda;
      32'H6052: READ <= 8'Hde;
      32'H6053: READ <= 8'He4;
      32'H6054: READ <= 8'He9;
      32'H6055: READ <= 8'Heb;
      32'H6056: READ <= 8'He6;
      32'H6057: READ <= 8'Heb;
      32'H6058: READ <= 8'He7;
      32'H6059: READ <= 8'Hac;
      32'H6060: READ <= 8'H1b;
      32'H6061: READ <= 8'H63;
      32'H6062: READ <= 8'H6e;
      32'H6063: READ <= 8'H5a;
      32'H6064: READ <= 8'H47;
      32'H6065: READ <= 8'H7a;
      32'H6066: READ <= 8'H78;
      32'H6067: READ <= 8'H97;
      32'H6068: READ <= 8'H9d;
      32'H6069: READ <= 8'Ha7;
      32'H6070: READ <= 8'H9d;
      32'H6071: READ <= 8'H89;
      32'H6072: READ <= 8'H77;
      32'H6073: READ <= 8'H73;
      32'H6074: READ <= 8'H75;
      32'H6075: READ <= 8'H76;
      32'H6076: READ <= 8'H77;
      32'H6077: READ <= 8'H78;
      32'H6078: READ <= 8'H79;
      32'H6079: READ <= 8'H7a;
      32'H6080: READ <= 8'H7b;
      32'H6081: READ <= 8'H7b;
      32'H6082: READ <= 8'H7c;
      32'H6083: READ <= 8'H7d;
      32'H6084: READ <= 8'H7d;
      32'H6085: READ <= 8'H7e;
      32'H6086: READ <= 8'H7f;
      32'H6087: READ <= 8'H80;
      32'H6088: READ <= 8'H81;
      32'H6089: READ <= 8'H82;
      32'H6090: READ <= 8'H83;
      32'H6091: READ <= 8'H84;
      32'H6092: READ <= 8'H85;
      32'H6093: READ <= 8'H86;
      32'H6094: READ <= 8'H87;
      32'H6095: READ <= 8'H87;
      32'H6096: READ <= 8'H87;
      32'H6097: READ <= 8'H88;
      32'H6098: READ <= 8'H89;
      32'H6099: READ <= 8'H8a;
      32'H6100: READ <= 8'H72;
      32'H6101: READ <= 8'H72;
      32'H6102: READ <= 8'H71;
      32'H6103: READ <= 8'H71;
      32'H6104: READ <= 8'H70;
      32'H6105: READ <= 8'H6f;
      32'H6106: READ <= 8'H6f;
      32'H6107: READ <= 8'H6e;
      32'H6108: READ <= 8'H6e;
      32'H6109: READ <= 8'H6e;
      32'H6110: READ <= 8'H6d;
      32'H6111: READ <= 8'H6c;
      32'H6112: READ <= 8'H6c;
      32'H6113: READ <= 8'H6b;
      32'H6114: READ <= 8'H6a;
      32'H6115: READ <= 8'H6a;
      32'H6116: READ <= 8'H6a;
      32'H6117: READ <= 8'H69;
      32'H6118: READ <= 8'H69;
      32'H6119: READ <= 8'H69;
      32'H6120: READ <= 8'H68;
      32'H6121: READ <= 8'H69;
      32'H6122: READ <= 8'H6a;
      32'H6123: READ <= 8'H6c;
      32'H6124: READ <= 8'H6e;
      32'H6125: READ <= 8'H70;
      32'H6126: READ <= 8'H74;
      32'H6127: READ <= 8'H79;
      32'H6128: READ <= 8'H7e;
      32'H6129: READ <= 8'H83;
      32'H6130: READ <= 8'H89;
      32'H6131: READ <= 8'H8d;
      32'H6132: READ <= 8'H90;
      32'H6133: READ <= 8'H96;
      32'H6134: READ <= 8'H88;
      32'H6135: READ <= 8'H77;
      32'H6136: READ <= 8'Hc3;
      32'H6137: READ <= 8'Hbd;
      32'H6138: READ <= 8'Ha1;
      32'H6139: READ <= 8'H81;
      32'H6140: READ <= 8'Hce;
      32'H6141: READ <= 8'Hd8;
      32'H6142: READ <= 8'Hd4;
      32'H6143: READ <= 8'Hd0;
      32'H6144: READ <= 8'Hce;
      32'H6145: READ <= 8'Hce;
      32'H6146: READ <= 8'Hcf;
      32'H6147: READ <= 8'Hcf;
      32'H6148: READ <= 8'Hcf;
      32'H6149: READ <= 8'Hd1;
      32'H6150: READ <= 8'Hd5;
      32'H6151: READ <= 8'Hd9;
      32'H6152: READ <= 8'Hdd;
      32'H6153: READ <= 8'He2;
      32'H6154: READ <= 8'He7;
      32'H6155: READ <= 8'He9;
      32'H6156: READ <= 8'He7;
      32'H6157: READ <= 8'Hec;
      32'H6158: READ <= 8'He0;
      32'H6159: READ <= 8'Hb2;
      32'H6160: READ <= 8'H23;
      32'H6161: READ <= 8'H66;
      32'H6162: READ <= 8'H4b;
      32'H6163: READ <= 8'H5c;
      32'H6164: READ <= 8'H54;
      32'H6165: READ <= 8'H83;
      32'H6166: READ <= 8'H8b;
      32'H6167: READ <= 8'H9d;
      32'H6168: READ <= 8'H95;
      32'H6169: READ <= 8'H90;
      32'H6170: READ <= 8'H90;
      32'H6171: READ <= 8'H76;
      32'H6172: READ <= 8'H72;
      32'H6173: READ <= 8'H74;
      32'H6174: READ <= 8'H75;
      32'H6175: READ <= 8'H76;
      32'H6176: READ <= 8'H76;
      32'H6177: READ <= 8'H78;
      32'H6178: READ <= 8'H79;
      32'H6179: READ <= 8'H7a;
      32'H6180: READ <= 8'H7a;
      32'H6181: READ <= 8'H7b;
      32'H6182: READ <= 8'H7b;
      32'H6183: READ <= 8'H7d;
      32'H6184: READ <= 8'H7d;
      32'H6185: READ <= 8'H7e;
      32'H6186: READ <= 8'H7f;
      32'H6187: READ <= 8'H80;
      32'H6188: READ <= 8'H80;
      32'H6189: READ <= 8'H81;
      32'H6190: READ <= 8'H83;
      32'H6191: READ <= 8'H84;
      32'H6192: READ <= 8'H85;
      32'H6193: READ <= 8'H86;
      32'H6194: READ <= 8'H87;
      32'H6195: READ <= 8'H88;
      32'H6196: READ <= 8'H87;
      32'H6197: READ <= 8'H88;
      32'H6198: READ <= 8'H88;
      32'H6199: READ <= 8'H89;
      32'H6200: READ <= 8'H72;
      32'H6201: READ <= 8'H71;
      32'H6202: READ <= 8'H72;
      32'H6203: READ <= 8'H71;
      32'H6204: READ <= 8'H70;
      32'H6205: READ <= 8'H70;
      32'H6206: READ <= 8'H6f;
      32'H6207: READ <= 8'H6f;
      32'H6208: READ <= 8'H6f;
      32'H6209: READ <= 8'H6e;
      32'H6210: READ <= 8'H6e;
      32'H6211: READ <= 8'H6d;
      32'H6212: READ <= 8'H6d;
      32'H6213: READ <= 8'H6c;
      32'H6214: READ <= 8'H6b;
      32'H6215: READ <= 8'H6a;
      32'H6216: READ <= 8'H6a;
      32'H6217: READ <= 8'H6a;
      32'H6218: READ <= 8'H6a;
      32'H6219: READ <= 8'H69;
      32'H6220: READ <= 8'H69;
      32'H6221: READ <= 8'H69;
      32'H6222: READ <= 8'H6a;
      32'H6223: READ <= 8'H6b;
      32'H6224: READ <= 8'H6b;
      32'H6225: READ <= 8'H6e;
      32'H6226: READ <= 8'H72;
      32'H6227: READ <= 8'H79;
      32'H6228: READ <= 8'H80;
      32'H6229: READ <= 8'H85;
      32'H6230: READ <= 8'H8b;
      32'H6231: READ <= 8'H8f;
      32'H6232: READ <= 8'H93;
      32'H6233: READ <= 8'H9c;
      32'H6234: READ <= 8'H74;
      32'H6235: READ <= 8'H94;
      32'H6236: READ <= 8'Hae;
      32'H6237: READ <= 8'Hb6;
      32'H6238: READ <= 8'Ha0;
      32'H6239: READ <= 8'H80;
      32'H6240: READ <= 8'Hc9;
      32'H6241: READ <= 8'Hd7;
      32'H6242: READ <= 8'Hd2;
      32'H6243: READ <= 8'Hd0;
      32'H6244: READ <= 8'Hce;
      32'H6245: READ <= 8'Hcf;
      32'H6246: READ <= 8'Hcf;
      32'H6247: READ <= 8'Hcf;
      32'H6248: READ <= 8'Hcf;
      32'H6249: READ <= 8'Hd1;
      32'H6250: READ <= 8'Hd4;
      32'H6251: READ <= 8'Hd8;
      32'H6252: READ <= 8'Hda;
      32'H6253: READ <= 8'Hde;
      32'H6254: READ <= 8'He2;
      32'H6255: READ <= 8'He5;
      32'H6256: READ <= 8'He5;
      32'H6257: READ <= 8'Hec;
      32'H6258: READ <= 8'Hd6;
      32'H6259: READ <= 8'H9b;
      32'H6260: READ <= 8'H62;
      32'H6261: READ <= 8'H7f;
      32'H6262: READ <= 8'H58;
      32'H6263: READ <= 8'H49;
      32'H6264: READ <= 8'H5a;
      32'H6265: READ <= 8'H91;
      32'H6266: READ <= 8'H8c;
      32'H6267: READ <= 8'H8f;
      32'H6268: READ <= 8'H9e;
      32'H6269: READ <= 8'H8f;
      32'H6270: READ <= 8'H76;
      32'H6271: READ <= 8'H71;
      32'H6272: READ <= 8'H71;
      32'H6273: READ <= 8'H73;
      32'H6274: READ <= 8'H74;
      32'H6275: READ <= 8'H76;
      32'H6276: READ <= 8'H77;
      32'H6277: READ <= 8'H78;
      32'H6278: READ <= 8'H79;
      32'H6279: READ <= 8'H7a;
      32'H6280: READ <= 8'H7a;
      32'H6281: READ <= 8'H7b;
      32'H6282: READ <= 8'H7c;
      32'H6283: READ <= 8'H7c;
      32'H6284: READ <= 8'H7d;
      32'H6285: READ <= 8'H7e;
      32'H6286: READ <= 8'H7f;
      32'H6287: READ <= 8'H80;
      32'H6288: READ <= 8'H80;
      32'H6289: READ <= 8'H82;
      32'H6290: READ <= 8'H83;
      32'H6291: READ <= 8'H84;
      32'H6292: READ <= 8'H85;
      32'H6293: READ <= 8'H86;
      32'H6294: READ <= 8'H87;
      32'H6295: READ <= 8'H87;
      32'H6296: READ <= 8'H87;
      32'H6297: READ <= 8'H88;
      32'H6298: READ <= 8'H88;
      32'H6299: READ <= 8'H89;
      32'H6300: READ <= 8'H72;
      32'H6301: READ <= 8'H72;
      32'H6302: READ <= 8'H71;
      32'H6303: READ <= 8'H70;
      32'H6304: READ <= 8'H70;
      32'H6305: READ <= 8'H70;
      32'H6306: READ <= 8'H70;
      32'H6307: READ <= 8'H6f;
      32'H6308: READ <= 8'H6f;
      32'H6309: READ <= 8'H6f;
      32'H6310: READ <= 8'H6e;
      32'H6311: READ <= 8'H6e;
      32'H6312: READ <= 8'H6d;
      32'H6313: READ <= 8'H6c;
      32'H6314: READ <= 8'H6c;
      32'H6315: READ <= 8'H6b;
      32'H6316: READ <= 8'H6a;
      32'H6317: READ <= 8'H6a;
      32'H6318: READ <= 8'H6a;
      32'H6319: READ <= 8'H6a;
      32'H6320: READ <= 8'H6a;
      32'H6321: READ <= 8'H6a;
      32'H6322: READ <= 8'H6a;
      32'H6323: READ <= 8'H6b;
      32'H6324: READ <= 8'H6b;
      32'H6325: READ <= 8'H6e;
      32'H6326: READ <= 8'H72;
      32'H6327: READ <= 8'H79;
      32'H6328: READ <= 8'H81;
      32'H6329: READ <= 8'H88;
      32'H6330: READ <= 8'H8e;
      32'H6331: READ <= 8'H92;
      32'H6332: READ <= 8'H96;
      32'H6333: READ <= 8'H9a;
      32'H6334: READ <= 8'H81;
      32'H6335: READ <= 8'H96;
      32'H6336: READ <= 8'Hc0;
      32'H6337: READ <= 8'Hcb;
      32'H6338: READ <= 8'Hae;
      32'H6339: READ <= 8'H8d;
      32'H6340: READ <= 8'Hc4;
      32'H6341: READ <= 8'Hd3;
      32'H6342: READ <= 8'Hd0;
      32'H6343: READ <= 8'Hcf;
      32'H6344: READ <= 8'Hcd;
      32'H6345: READ <= 8'Hcf;
      32'H6346: READ <= 8'Hcf;
      32'H6347: READ <= 8'Hce;
      32'H6348: READ <= 8'Hce;
      32'H6349: READ <= 8'Hd0;
      32'H6350: READ <= 8'Hd3;
      32'H6351: READ <= 8'Hd6;
      32'H6352: READ <= 8'Hd8;
      32'H6353: READ <= 8'Hda;
      32'H6354: READ <= 8'Hdb;
      32'H6355: READ <= 8'Hdb;
      32'H6356: READ <= 8'He3;
      32'H6357: READ <= 8'He8;
      32'H6358: READ <= 8'Hd3;
      32'H6359: READ <= 8'H61;
      32'H6360: READ <= 8'H77;
      32'H6361: READ <= 8'H93;
      32'H6362: READ <= 8'H57;
      32'H6363: READ <= 8'H53;
      32'H6364: READ <= 8'H80;
      32'H6365: READ <= 8'H94;
      32'H6366: READ <= 8'H98;
      32'H6367: READ <= 8'H8f;
      32'H6368: READ <= 8'H7d;
      32'H6369: READ <= 8'H73;
      32'H6370: READ <= 8'H70;
      32'H6371: READ <= 8'H71;
      32'H6372: READ <= 8'H71;
      32'H6373: READ <= 8'H72;
      32'H6374: READ <= 8'H74;
      32'H6375: READ <= 8'H75;
      32'H6376: READ <= 8'H76;
      32'H6377: READ <= 8'H78;
      32'H6378: READ <= 8'H78;
      32'H6379: READ <= 8'H7a;
      32'H6380: READ <= 8'H7a;
      32'H6381: READ <= 8'H7b;
      32'H6382: READ <= 8'H7c;
      32'H6383: READ <= 8'H7c;
      32'H6384: READ <= 8'H7d;
      32'H6385: READ <= 8'H7e;
      32'H6386: READ <= 8'H7e;
      32'H6387: READ <= 8'H80;
      32'H6388: READ <= 8'H80;
      32'H6389: READ <= 8'H82;
      32'H6390: READ <= 8'H83;
      32'H6391: READ <= 8'H84;
      32'H6392: READ <= 8'H84;
      32'H6393: READ <= 8'H85;
      32'H6394: READ <= 8'H86;
      32'H6395: READ <= 8'H87;
      32'H6396: READ <= 8'H87;
      32'H6397: READ <= 8'H88;
      32'H6398: READ <= 8'H88;
      32'H6399: READ <= 8'H88;
      32'H6400: READ <= 8'H72;
      32'H6401: READ <= 8'H71;
      32'H6402: READ <= 8'H72;
      32'H6403: READ <= 8'H71;
      32'H6404: READ <= 8'H71;
      32'H6405: READ <= 8'H70;
      32'H6406: READ <= 8'H70;
      32'H6407: READ <= 8'H70;
      32'H6408: READ <= 8'H70;
      32'H6409: READ <= 8'H6f;
      32'H6410: READ <= 8'H6e;
      32'H6411: READ <= 8'H6e;
      32'H6412: READ <= 8'H6d;
      32'H6413: READ <= 8'H6d;
      32'H6414: READ <= 8'H6c;
      32'H6415: READ <= 8'H6c;
      32'H6416: READ <= 8'H6b;
      32'H6417: READ <= 8'H6b;
      32'H6418: READ <= 8'H6b;
      32'H6419: READ <= 8'H6b;
      32'H6420: READ <= 8'H6b;
      32'H6421: READ <= 8'H6b;
      32'H6422: READ <= 8'H6b;
      32'H6423: READ <= 8'H6b;
      32'H6424: READ <= 8'H6b;
      32'H6425: READ <= 8'H6e;
      32'H6426: READ <= 8'H73;
      32'H6427: READ <= 8'H7a;
      32'H6428: READ <= 8'H82;
      32'H6429: READ <= 8'H8a;
      32'H6430: READ <= 8'H90;
      32'H6431: READ <= 8'H94;
      32'H6432: READ <= 8'H99;
      32'H6433: READ <= 8'H92;
      32'H6434: READ <= 8'H85;
      32'H6435: READ <= 8'Hab;
      32'H6436: READ <= 8'Hca;
      32'H6437: READ <= 8'Hdb;
      32'H6438: READ <= 8'Hc3;
      32'H6439: READ <= 8'Ha3;
      32'H6440: READ <= 8'Hbc;
      32'H6441: READ <= 8'Hcd;
      32'H6442: READ <= 8'Hce;
      32'H6443: READ <= 8'Hcf;
      32'H6444: READ <= 8'Hcd;
      32'H6445: READ <= 8'Hce;
      32'H6446: READ <= 8'Hcf;
      32'H6447: READ <= 8'Hcd;
      32'H6448: READ <= 8'Hcd;
      32'H6449: READ <= 8'Hce;
      32'H6450: READ <= 8'Hd1;
      32'H6451: READ <= 8'Hd3;
      32'H6452: READ <= 8'Hd6;
      32'H6453: READ <= 8'Hd8;
      32'H6454: READ <= 8'Hd6;
      32'H6455: READ <= 8'Hcc;
      32'H6456: READ <= 8'Hde;
      32'H6457: READ <= 8'Hd6;
      32'H6458: READ <= 8'Haa;
      32'H6459: READ <= 8'H5a;
      32'H6460: READ <= 8'Ha4;
      32'H6461: READ <= 8'H9f;
      32'H6462: READ <= 8'H8e;
      32'H6463: READ <= 8'H91;
      32'H6464: READ <= 8'Had;
      32'H6465: READ <= 8'H91;
      32'H6466: READ <= 8'H94;
      32'H6467: READ <= 8'H7a;
      32'H6468: READ <= 8'H78;
      32'H6469: READ <= 8'H73;
      32'H6470: READ <= 8'H71;
      32'H6471: READ <= 8'H71;
      32'H6472: READ <= 8'H72;
      32'H6473: READ <= 8'H73;
      32'H6474: READ <= 8'H74;
      32'H6475: READ <= 8'H75;
      32'H6476: READ <= 8'H76;
      32'H6477: READ <= 8'H77;
      32'H6478: READ <= 8'H78;
      32'H6479: READ <= 8'H79;
      32'H6480: READ <= 8'H7b;
      32'H6481: READ <= 8'H7b;
      32'H6482: READ <= 8'H7c;
      32'H6483: READ <= 8'H7c;
      32'H6484: READ <= 8'H7d;
      32'H6485: READ <= 8'H7d;
      32'H6486: READ <= 8'H7e;
      32'H6487: READ <= 8'H7f;
      32'H6488: READ <= 8'H80;
      32'H6489: READ <= 8'H81;
      32'H6490: READ <= 8'H83;
      32'H6491: READ <= 8'H84;
      32'H6492: READ <= 8'H84;
      32'H6493: READ <= 8'H85;
      32'H6494: READ <= 8'H86;
      32'H6495: READ <= 8'H86;
      32'H6496: READ <= 8'H87;
      32'H6497: READ <= 8'H88;
      32'H6498: READ <= 8'H88;
      32'H6499: READ <= 8'H88;
      32'H6500: READ <= 8'H73;
      32'H6501: READ <= 8'H72;
      32'H6502: READ <= 8'H72;
      32'H6503: READ <= 8'H71;
      32'H6504: READ <= 8'H71;
      32'H6505: READ <= 8'H70;
      32'H6506: READ <= 8'H70;
      32'H6507: READ <= 8'H70;
      32'H6508: READ <= 8'H70;
      32'H6509: READ <= 8'H6f;
      32'H6510: READ <= 8'H6f;
      32'H6511: READ <= 8'H6f;
      32'H6512: READ <= 8'H6e;
      32'H6513: READ <= 8'H6d;
      32'H6514: READ <= 8'H6d;
      32'H6515: READ <= 8'H6d;
      32'H6516: READ <= 8'H6c;
      32'H6517: READ <= 8'H6c;
      32'H6518: READ <= 8'H6c;
      32'H6519: READ <= 8'H6b;
      32'H6520: READ <= 8'H6c;
      32'H6521: READ <= 8'H6b;
      32'H6522: READ <= 8'H6c;
      32'H6523: READ <= 8'H6c;
      32'H6524: READ <= 8'H6c;
      32'H6525: READ <= 8'H70;
      32'H6526: READ <= 8'H75;
      32'H6527: READ <= 8'H7c;
      32'H6528: READ <= 8'H85;
      32'H6529: READ <= 8'H8c;
      32'H6530: READ <= 8'H92;
      32'H6531: READ <= 8'H97;
      32'H6532: READ <= 8'H99;
      32'H6533: READ <= 8'H7f;
      32'H6534: READ <= 8'H9a;
      32'H6535: READ <= 8'Hd1;
      32'H6536: READ <= 8'Hd0;
      32'H6537: READ <= 8'Hdb;
      32'H6538: READ <= 8'Hcd;
      32'H6539: READ <= 8'Hb9;
      32'H6540: READ <= 8'Hbc;
      32'H6541: READ <= 8'Hc8;
      32'H6542: READ <= 8'Hcd;
      32'H6543: READ <= 8'Hd0;
      32'H6544: READ <= 8'Hce;
      32'H6545: READ <= 8'Hce;
      32'H6546: READ <= 8'Hcf;
      32'H6547: READ <= 8'Hcd;
      32'H6548: READ <= 8'Hcc;
      32'H6549: READ <= 8'Hcc;
      32'H6550: READ <= 8'Hce;
      32'H6551: READ <= 8'Hd0;
      32'H6552: READ <= 8'Hd2;
      32'H6553: READ <= 8'Hd5;
      32'H6554: READ <= 8'Hd8;
      32'H6555: READ <= 8'Hcf;
      32'H6556: READ <= 8'Hdd;
      32'H6557: READ <= 8'Hb5;
      32'H6558: READ <= 8'H68;
      32'H6559: READ <= 8'Ha2;
      32'H6560: READ <= 8'Hb5;
      32'H6561: READ <= 8'Ha9;
      32'H6562: READ <= 8'H9b;
      32'H6563: READ <= 8'H98;
      32'H6564: READ <= 8'H87;
      32'H6565: READ <= 8'H82;
      32'H6566: READ <= 8'H7f;
      32'H6567: READ <= 8'H7d;
      32'H6568: READ <= 8'H78;
      32'H6569: READ <= 8'H75;
      32'H6570: READ <= 8'H72;
      32'H6571: READ <= 8'H71;
      32'H6572: READ <= 8'H71;
      32'H6573: READ <= 8'H72;
      32'H6574: READ <= 8'H74;
      32'H6575: READ <= 8'H75;
      32'H6576: READ <= 8'H76;
      32'H6577: READ <= 8'H78;
      32'H6578: READ <= 8'H79;
      32'H6579: READ <= 8'H7a;
      32'H6580: READ <= 8'H7a;
      32'H6581: READ <= 8'H7a;
      32'H6582: READ <= 8'H7b;
      32'H6583: READ <= 8'H7c;
      32'H6584: READ <= 8'H7d;
      32'H6585: READ <= 8'H7d;
      32'H6586: READ <= 8'H7e;
      32'H6587: READ <= 8'H80;
      32'H6588: READ <= 8'H80;
      32'H6589: READ <= 8'H82;
      32'H6590: READ <= 8'H82;
      32'H6591: READ <= 8'H83;
      32'H6592: READ <= 8'H85;
      32'H6593: READ <= 8'H85;
      32'H6594: READ <= 8'H86;
      32'H6595: READ <= 8'H86;
      32'H6596: READ <= 8'H86;
      32'H6597: READ <= 8'H88;
      32'H6598: READ <= 8'H88;
      32'H6599: READ <= 8'H88;
      32'H6600: READ <= 8'H73;
      32'H6601: READ <= 8'H73;
      32'H6602: READ <= 8'H73;
      32'H6603: READ <= 8'H72;
      32'H6604: READ <= 8'H72;
      32'H6605: READ <= 8'H71;
      32'H6606: READ <= 8'H70;
      32'H6607: READ <= 8'H70;
      32'H6608: READ <= 8'H70;
      32'H6609: READ <= 8'H70;
      32'H6610: READ <= 8'H70;
      32'H6611: READ <= 8'H6f;
      32'H6612: READ <= 8'H6f;
      32'H6613: READ <= 8'H6f;
      32'H6614: READ <= 8'H6e;
      32'H6615: READ <= 8'H6d;
      32'H6616: READ <= 8'H6c;
      32'H6617: READ <= 8'H6d;
      32'H6618: READ <= 8'H6d;
      32'H6619: READ <= 8'H6c;
      32'H6620: READ <= 8'H6c;
      32'H6621: READ <= 8'H6c;
      32'H6622: READ <= 8'H6c;
      32'H6623: READ <= 8'H6c;
      32'H6624: READ <= 8'H6e;
      32'H6625: READ <= 8'H71;
      32'H6626: READ <= 8'H77;
      32'H6627: READ <= 8'H7e;
      32'H6628: READ <= 8'H87;
      32'H6629: READ <= 8'H8e;
      32'H6630: READ <= 8'H95;
      32'H6631: READ <= 8'H98;
      32'H6632: READ <= 8'H98;
      32'H6633: READ <= 8'H80;
      32'H6634: READ <= 8'Ha0;
      32'H6635: READ <= 8'Hdf;
      32'H6636: READ <= 8'Hd9;
      32'H6637: READ <= 8'Hd9;
      32'H6638: READ <= 8'Hd4;
      32'H6639: READ <= 8'Hc9;
      32'H6640: READ <= 8'Hc4;
      32'H6641: READ <= 8'Hc7;
      32'H6642: READ <= 8'Hcf;
      32'H6643: READ <= 8'Hd2;
      32'H6644: READ <= 8'Hd0;
      32'H6645: READ <= 8'Hcf;
      32'H6646: READ <= 8'Hcf;
      32'H6647: READ <= 8'Hce;
      32'H6648: READ <= 8'Hcd;
      32'H6649: READ <= 8'Hcc;
      32'H6650: READ <= 8'Hcc;
      32'H6651: READ <= 8'Hcc;
      32'H6652: READ <= 8'Hcd;
      32'H6653: READ <= 8'Hd0;
      32'H6654: READ <= 8'Hda;
      32'H6655: READ <= 8'Hdc;
      32'H6656: READ <= 8'Hcd;
      32'H6657: READ <= 8'Ha1;
      32'H6658: READ <= 8'H91;
      32'H6659: READ <= 8'Hc0;
      32'H6660: READ <= 8'Hba;
      32'H6661: READ <= 8'Hb1;
      32'H6662: READ <= 8'Ha4;
      32'H6663: READ <= 8'H97;
      32'H6664: READ <= 8'H8f;
      32'H6665: READ <= 8'H89;
      32'H6666: READ <= 8'H84;
      32'H6667: READ <= 8'H7f;
      32'H6668: READ <= 8'H7c;
      32'H6669: READ <= 8'H78;
      32'H6670: READ <= 8'H75;
      32'H6671: READ <= 8'H72;
      32'H6672: READ <= 8'H72;
      32'H6673: READ <= 8'H72;
      32'H6674: READ <= 8'H73;
      32'H6675: READ <= 8'H75;
      32'H6676: READ <= 8'H76;
      32'H6677: READ <= 8'H77;
      32'H6678: READ <= 8'H78;
      32'H6679: READ <= 8'H79;
      32'H6680: READ <= 8'H7a;
      32'H6681: READ <= 8'H7a;
      32'H6682: READ <= 8'H7c;
      32'H6683: READ <= 8'H7c;
      32'H6684: READ <= 8'H7d;
      32'H6685: READ <= 8'H7e;
      32'H6686: READ <= 8'H7f;
      32'H6687: READ <= 8'H7f;
      32'H6688: READ <= 8'H81;
      32'H6689: READ <= 8'H81;
      32'H6690: READ <= 8'H82;
      32'H6691: READ <= 8'H83;
      32'H6692: READ <= 8'H84;
      32'H6693: READ <= 8'H85;
      32'H6694: READ <= 8'H86;
      32'H6695: READ <= 8'H86;
      32'H6696: READ <= 8'H86;
      32'H6697: READ <= 8'H87;
      32'H6698: READ <= 8'H88;
      32'H6699: READ <= 8'H88;
      32'H6700: READ <= 8'H73;
      32'H6701: READ <= 8'H73;
      32'H6702: READ <= 8'H73;
      32'H6703: READ <= 8'H73;
      32'H6704: READ <= 8'H72;
      32'H6705: READ <= 8'H71;
      32'H6706: READ <= 8'H70;
      32'H6707: READ <= 8'H70;
      32'H6708: READ <= 8'H70;
      32'H6709: READ <= 8'H70;
      32'H6710: READ <= 8'H70;
      32'H6711: READ <= 8'H70;
      32'H6712: READ <= 8'H6f;
      32'H6713: READ <= 8'H6f;
      32'H6714: READ <= 8'H6e;
      32'H6715: READ <= 8'H6d;
      32'H6716: READ <= 8'H6d;
      32'H6717: READ <= 8'H6e;
      32'H6718: READ <= 8'H6d;
      32'H6719: READ <= 8'H6d;
      32'H6720: READ <= 8'H6e;
      32'H6721: READ <= 8'H6d;
      32'H6722: READ <= 8'H6d;
      32'H6723: READ <= 8'H6d;
      32'H6724: READ <= 8'H6e;
      32'H6725: READ <= 8'H73;
      32'H6726: READ <= 8'H79;
      32'H6727: READ <= 8'H7f;
      32'H6728: READ <= 8'H89;
      32'H6729: READ <= 8'H90;
      32'H6730: READ <= 8'H96;
      32'H6731: READ <= 8'H98;
      32'H6732: READ <= 8'H9c;
      32'H6733: READ <= 8'H7f;
      32'H6734: READ <= 8'Ha9;
      32'H6735: READ <= 8'He1;
      32'H6736: READ <= 8'He1;
      32'H6737: READ <= 8'Hdd;
      32'H6738: READ <= 8'Hd8;
      32'H6739: READ <= 8'Hd4;
      32'H6740: READ <= 8'Hce;
      32'H6741: READ <= 8'Hcd;
      32'H6742: READ <= 8'Hd1;
      32'H6743: READ <= 8'Hd4;
      32'H6744: READ <= 8'Hd3;
      32'H6745: READ <= 8'Hd1;
      32'H6746: READ <= 8'Hd0;
      32'H6747: READ <= 8'Hd0;
      32'H6748: READ <= 8'Hce;
      32'H6749: READ <= 8'Hcd;
      32'H6750: READ <= 8'Hcb;
      32'H6751: READ <= 8'Hca;
      32'H6752: READ <= 8'Hc8;
      32'H6753: READ <= 8'Hca;
      32'H6754: READ <= 8'Hd7;
      32'H6755: READ <= 8'He2;
      32'H6756: READ <= 8'Hc7;
      32'H6757: READ <= 8'H91;
      32'H6758: READ <= 8'Haf;
      32'H6759: READ <= 8'Hc5;
      32'H6760: READ <= 8'Hbf;
      32'H6761: READ <= 8'Hb7;
      32'H6762: READ <= 8'Hab;
      32'H6763: READ <= 8'H9d;
      32'H6764: READ <= 8'H94;
      32'H6765: READ <= 8'H8c;
      32'H6766: READ <= 8'H87;
      32'H6767: READ <= 8'H82;
      32'H6768: READ <= 8'H7f;
      32'H6769: READ <= 8'H7a;
      32'H6770: READ <= 8'H77;
      32'H6771: READ <= 8'H74;
      32'H6772: READ <= 8'H73;
      32'H6773: READ <= 8'H73;
      32'H6774: READ <= 8'H73;
      32'H6775: READ <= 8'H74;
      32'H6776: READ <= 8'H76;
      32'H6777: READ <= 8'H76;
      32'H6778: READ <= 8'H78;
      32'H6779: READ <= 8'H78;
      32'H6780: READ <= 8'H7a;
      32'H6781: READ <= 8'H7a;
      32'H6782: READ <= 8'H7b;
      32'H6783: READ <= 8'H7c;
      32'H6784: READ <= 8'H7d;
      32'H6785: READ <= 8'H7e;
      32'H6786: READ <= 8'H7f;
      32'H6787: READ <= 8'H7f;
      32'H6788: READ <= 8'H81;
      32'H6789: READ <= 8'H81;
      32'H6790: READ <= 8'H82;
      32'H6791: READ <= 8'H83;
      32'H6792: READ <= 8'H84;
      32'H6793: READ <= 8'H84;
      32'H6794: READ <= 8'H85;
      32'H6795: READ <= 8'H85;
      32'H6796: READ <= 8'H86;
      32'H6797: READ <= 8'H87;
      32'H6798: READ <= 8'H88;
      32'H6799: READ <= 8'H88;
      32'H6800: READ <= 8'H74;
      32'H6801: READ <= 8'H74;
      32'H6802: READ <= 8'H74;
      32'H6803: READ <= 8'H73;
      32'H6804: READ <= 8'H72;
      32'H6805: READ <= 8'H72;
      32'H6806: READ <= 8'H71;
      32'H6807: READ <= 8'H71;
      32'H6808: READ <= 8'H70;
      32'H6809: READ <= 8'H70;
      32'H6810: READ <= 8'H70;
      32'H6811: READ <= 8'H70;
      32'H6812: READ <= 8'H70;
      32'H6813: READ <= 8'H70;
      32'H6814: READ <= 8'H6f;
      32'H6815: READ <= 8'H6e;
      32'H6816: READ <= 8'H6e;
      32'H6817: READ <= 8'H6e;
      32'H6818: READ <= 8'H6e;
      32'H6819: READ <= 8'H6e;
      32'H6820: READ <= 8'H6d;
      32'H6821: READ <= 8'H6d;
      32'H6822: READ <= 8'H6d;
      32'H6823: READ <= 8'H6d;
      32'H6824: READ <= 8'H6e;
      32'H6825: READ <= 8'H74;
      32'H6826: READ <= 8'H7a;
      32'H6827: READ <= 8'H80;
      32'H6828: READ <= 8'H89;
      32'H6829: READ <= 8'H91;
      32'H6830: READ <= 8'H97;
      32'H6831: READ <= 8'H98;
      32'H6832: READ <= 8'Ha8;
      32'H6833: READ <= 8'H8e;
      32'H6834: READ <= 8'Hcf;
      32'H6835: READ <= 8'He5;
      32'H6836: READ <= 8'He6;
      32'H6837: READ <= 8'He4;
      32'H6838: READ <= 8'Hdd;
      32'H6839: READ <= 8'Hda;
      32'H6840: READ <= 8'Hd8;
      32'H6841: READ <= 8'Hd6;
      32'H6842: READ <= 8'Hd6;
      32'H6843: READ <= 8'Hd5;
      32'H6844: READ <= 8'Hd5;
      32'H6845: READ <= 8'Hd4;
      32'H6846: READ <= 8'Hd3;
      32'H6847: READ <= 8'Hd3;
      32'H6848: READ <= 8'Hd1;
      32'H6849: READ <= 8'Hcf;
      32'H6850: READ <= 8'Hcd;
      32'H6851: READ <= 8'Hcb;
      32'H6852: READ <= 8'Hc6;
      32'H6853: READ <= 8'Hc4;
      32'H6854: READ <= 8'Hce;
      32'H6855: READ <= 8'Hdc;
      32'H6856: READ <= 8'Hce;
      32'H6857: READ <= 8'H8b;
      32'H6858: READ <= 8'Hc8;
      32'H6859: READ <= 8'Hc9;
      32'H6860: READ <= 8'Hc3;
      32'H6861: READ <= 8'Hbb;
      32'H6862: READ <= 8'Hb0;
      32'H6863: READ <= 8'Ha3;
      32'H6864: READ <= 8'H98;
      32'H6865: READ <= 8'H91;
      32'H6866: READ <= 8'H8a;
      32'H6867: READ <= 8'H85;
      32'H6868: READ <= 8'H81;
      32'H6869: READ <= 8'H7d;
      32'H6870: READ <= 8'H79;
      32'H6871: READ <= 8'H77;
      32'H6872: READ <= 8'H74;
      32'H6873: READ <= 8'H73;
      32'H6874: READ <= 8'H73;
      32'H6875: READ <= 8'H75;
      32'H6876: READ <= 8'H76;
      32'H6877: READ <= 8'H76;
      32'H6878: READ <= 8'H78;
      32'H6879: READ <= 8'H79;
      32'H6880: READ <= 8'H79;
      32'H6881: READ <= 8'H7a;
      32'H6882: READ <= 8'H7b;
      32'H6883: READ <= 8'H7c;
      32'H6884: READ <= 8'H7d;
      32'H6885: READ <= 8'H7d;
      32'H6886: READ <= 8'H7f;
      32'H6887: READ <= 8'H80;
      32'H6888: READ <= 8'H81;
      32'H6889: READ <= 8'H81;
      32'H6890: READ <= 8'H82;
      32'H6891: READ <= 8'H83;
      32'H6892: READ <= 8'H84;
      32'H6893: READ <= 8'H84;
      32'H6894: READ <= 8'H85;
      32'H6895: READ <= 8'H86;
      32'H6896: READ <= 8'H86;
      32'H6897: READ <= 8'H87;
      32'H6898: READ <= 8'H88;
      32'H6899: READ <= 8'H88;
      32'H6900: READ <= 8'H74;
      32'H6901: READ <= 8'H74;
      32'H6902: READ <= 8'H74;
      32'H6903: READ <= 8'H74;
      32'H6904: READ <= 8'H74;
      32'H6905: READ <= 8'H73;
      32'H6906: READ <= 8'H72;
      32'H6907: READ <= 8'H72;
      32'H6908: READ <= 8'H72;
      32'H6909: READ <= 8'H71;
      32'H6910: READ <= 8'H71;
      32'H6911: READ <= 8'H70;
      32'H6912: READ <= 8'H70;
      32'H6913: READ <= 8'H70;
      32'H6914: READ <= 8'H6f;
      32'H6915: READ <= 8'H6f;
      32'H6916: READ <= 8'H6f;
      32'H6917: READ <= 8'H6f;
      32'H6918: READ <= 8'H6e;
      32'H6919: READ <= 8'H6e;
      32'H6920: READ <= 8'H6e;
      32'H6921: READ <= 8'H6e;
      32'H6922: READ <= 8'H6d;
      32'H6923: READ <= 8'H6e;
      32'H6924: READ <= 8'H6f;
      32'H6925: READ <= 8'H74;
      32'H6926: READ <= 8'H7b;
      32'H6927: READ <= 8'H82;
      32'H6928: READ <= 8'H8a;
      32'H6929: READ <= 8'H92;
      32'H6930: READ <= 8'H98;
      32'H6931: READ <= 8'H9b;
      32'H6932: READ <= 8'Ha3;
      32'H6933: READ <= 8'Hae;
      32'H6934: READ <= 8'Hc7;
      32'H6935: READ <= 8'Hde;
      32'H6936: READ <= 8'He4;
      32'H6937: READ <= 8'He4;
      32'H6938: READ <= 8'Hdf;
      32'H6939: READ <= 8'Hdd;
      32'H6940: READ <= 8'Hdb;
      32'H6941: READ <= 8'Hda;
      32'H6942: READ <= 8'Hd8;
      32'H6943: READ <= 8'Hd5;
      32'H6944: READ <= 8'Hd4;
      32'H6945: READ <= 8'Hd4;
      32'H6946: READ <= 8'Hd4;
      32'H6947: READ <= 8'Hd4;
      32'H6948: READ <= 8'Hd1;
      32'H6949: READ <= 8'Hce;
      32'H6950: READ <= 8'Hcc;
      32'H6951: READ <= 8'Hca;
      32'H6952: READ <= 8'Hc7;
      32'H6953: READ <= 8'Hc5;
      32'H6954: READ <= 8'Hcc;
      32'H6955: READ <= 8'Hdc;
      32'H6956: READ <= 8'Ha3;
      32'H6957: READ <= 8'Ha8;
      32'H6958: READ <= 8'Hd3;
      32'H6959: READ <= 8'Hcd;
      32'H6960: READ <= 8'Hc6;
      32'H6961: READ <= 8'Hbf;
      32'H6962: READ <= 8'Hb5;
      32'H6963: READ <= 8'Ha9;
      32'H6964: READ <= 8'H9c;
      32'H6965: READ <= 8'H94;
      32'H6966: READ <= 8'H8e;
      32'H6967: READ <= 8'H88;
      32'H6968: READ <= 8'H84;
      32'H6969: READ <= 8'H80;
      32'H6970: READ <= 8'H7b;
      32'H6971: READ <= 8'H78;
      32'H6972: READ <= 8'H76;
      32'H6973: READ <= 8'H73;
      32'H6974: READ <= 8'H73;
      32'H6975: READ <= 8'H74;
      32'H6976: READ <= 8'H75;
      32'H6977: READ <= 8'H76;
      32'H6978: READ <= 8'H77;
      32'H6979: READ <= 8'H78;
      32'H6980: READ <= 8'H79;
      32'H6981: READ <= 8'H7a;
      32'H6982: READ <= 8'H7b;
      32'H6983: READ <= 8'H7c;
      32'H6984: READ <= 8'H7d;
      32'H6985: READ <= 8'H7d;
      32'H6986: READ <= 8'H7f;
      32'H6987: READ <= 8'H7f;
      32'H6988: READ <= 8'H80;
      32'H6989: READ <= 8'H81;
      32'H6990: READ <= 8'H82;
      32'H6991: READ <= 8'H82;
      32'H6992: READ <= 8'H83;
      32'H6993: READ <= 8'H84;
      32'H6994: READ <= 8'H85;
      32'H6995: READ <= 8'H86;
      32'H6996: READ <= 8'H86;
      32'H6997: READ <= 8'H87;
      32'H6998: READ <= 8'H88;
      32'H6999: READ <= 8'H88;
      32'H7000: READ <= 8'H74;
      32'H7001: READ <= 8'H74;
      32'H7002: READ <= 8'H74;
      32'H7003: READ <= 8'H74;
      32'H7004: READ <= 8'H74;
      32'H7005: READ <= 8'H74;
      32'H7006: READ <= 8'H73;
      32'H7007: READ <= 8'H73;
      32'H7008: READ <= 8'H73;
      32'H7009: READ <= 8'H71;
      32'H7010: READ <= 8'H72;
      32'H7011: READ <= 8'H71;
      32'H7012: READ <= 8'H71;
      32'H7013: READ <= 8'H71;
      32'H7014: READ <= 8'H70;
      32'H7015: READ <= 8'H6f;
      32'H7016: READ <= 8'H6f;
      32'H7017: READ <= 8'H6f;
      32'H7018: READ <= 8'H6f;
      32'H7019: READ <= 8'H6f;
      32'H7020: READ <= 8'H6e;
      32'H7021: READ <= 8'H6e;
      32'H7022: READ <= 8'H6e;
      32'H7023: READ <= 8'H6e;
      32'H7024: READ <= 8'H70;
      32'H7025: READ <= 8'H75;
      32'H7026: READ <= 8'H7b;
      32'H7027: READ <= 8'H84;
      32'H7028: READ <= 8'H8b;
      32'H7029: READ <= 8'H92;
      32'H7030: READ <= 8'H99;
      32'H7031: READ <= 8'H9f;
      32'H7032: READ <= 8'H9f;
      32'H7033: READ <= 8'Hb9;
      32'H7034: READ <= 8'Hb8;
      32'H7035: READ <= 8'Hcd;
      32'H7036: READ <= 8'Hdb;
      32'H7037: READ <= 8'Hdf;
      32'H7038: READ <= 8'Hde;
      32'H7039: READ <= 8'Hdc;
      32'H7040: READ <= 8'Hdc;
      32'H7041: READ <= 8'Hdc;
      32'H7042: READ <= 8'Hda;
      32'H7043: READ <= 8'Hd6;
      32'H7044: READ <= 8'Hd4;
      32'H7045: READ <= 8'Hd4;
      32'H7046: READ <= 8'Hd3;
      32'H7047: READ <= 8'Hd2;
      32'H7048: READ <= 8'Hd0;
      32'H7049: READ <= 8'Hce;
      32'H7050: READ <= 8'Hcd;
      32'H7051: READ <= 8'Hca;
      32'H7052: READ <= 8'Hc7;
      32'H7053: READ <= 8'Hc8;
      32'H7054: READ <= 8'Hce;
      32'H7055: READ <= 8'Hbf;
      32'H7056: READ <= 8'Haa;
      32'H7057: READ <= 8'Hcd;
      32'H7058: READ <= 8'Hd5;
      32'H7059: READ <= 8'Hce;
      32'H7060: READ <= 8'Hca;
      32'H7061: READ <= 8'Hc3;
      32'H7062: READ <= 8'Hb9;
      32'H7063: READ <= 8'Had;
      32'H7064: READ <= 8'Ha0;
      32'H7065: READ <= 8'H97;
      32'H7066: READ <= 8'H91;
      32'H7067: READ <= 8'H8b;
      32'H7068: READ <= 8'H86;
      32'H7069: READ <= 8'H82;
      32'H7070: READ <= 8'H7e;
      32'H7071: READ <= 8'H7a;
      32'H7072: READ <= 8'H78;
      32'H7073: READ <= 8'H75;
      32'H7074: READ <= 8'H74;
      32'H7075: READ <= 8'H74;
      32'H7076: READ <= 8'H75;
      32'H7077: READ <= 8'H76;
      32'H7078: READ <= 8'H77;
      32'H7079: READ <= 8'H78;
      32'H7080: READ <= 8'H79;
      32'H7081: READ <= 8'H7a;
      32'H7082: READ <= 8'H7b;
      32'H7083: READ <= 8'H7c;
      32'H7084: READ <= 8'H7d;
      32'H7085: READ <= 8'H7d;
      32'H7086: READ <= 8'H7e;
      32'H7087: READ <= 8'H7f;
      32'H7088: READ <= 8'H7f;
      32'H7089: READ <= 8'H81;
      32'H7090: READ <= 8'H81;
      32'H7091: READ <= 8'H82;
      32'H7092: READ <= 8'H84;
      32'H7093: READ <= 8'H84;
      32'H7094: READ <= 8'H85;
      32'H7095: READ <= 8'H86;
      32'H7096: READ <= 8'H86;
      32'H7097: READ <= 8'H87;
      32'H7098: READ <= 8'H87;
      32'H7099: READ <= 8'H87;
      32'H7100: READ <= 8'H75;
      32'H7101: READ <= 8'H75;
      32'H7102: READ <= 8'H75;
      32'H7103: READ <= 8'H75;
      32'H7104: READ <= 8'H75;
      32'H7105: READ <= 8'H75;
      32'H7106: READ <= 8'H74;
      32'H7107: READ <= 8'H74;
      32'H7108: READ <= 8'H73;
      32'H7109: READ <= 8'H73;
      32'H7110: READ <= 8'H73;
      32'H7111: READ <= 8'H71;
      32'H7112: READ <= 8'H71;
      32'H7113: READ <= 8'H71;
      32'H7114: READ <= 8'H70;
      32'H7115: READ <= 8'H70;
      32'H7116: READ <= 8'H70;
      32'H7117: READ <= 8'H6f;
      32'H7118: READ <= 8'H6f;
      32'H7119: READ <= 8'H6f;
      32'H7120: READ <= 8'H6f;
      32'H7121: READ <= 8'H6e;
      32'H7122: READ <= 8'H6f;
      32'H7123: READ <= 8'H6f;
      32'H7124: READ <= 8'H71;
      32'H7125: READ <= 8'H76;
      32'H7126: READ <= 8'H7c;
      32'H7127: READ <= 8'H85;
      32'H7128: READ <= 8'H8e;
      32'H7129: READ <= 8'H94;
      32'H7130: READ <= 8'H9d;
      32'H7131: READ <= 8'Ha3;
      32'H7132: READ <= 8'Hb5;
      32'H7133: READ <= 8'Hba;
      32'H7134: READ <= 8'Hb7;
      32'H7135: READ <= 8'Hc1;
      32'H7136: READ <= 8'Hd0;
      32'H7137: READ <= 8'Hd9;
      32'H7138: READ <= 8'Hda;
      32'H7139: READ <= 8'Hdb;
      32'H7140: READ <= 8'Hdc;
      32'H7141: READ <= 8'Hdc;
      32'H7142: READ <= 8'Hdd;
      32'H7143: READ <= 8'Hd8;
      32'H7144: READ <= 8'Hd6;
      32'H7145: READ <= 8'Hd6;
      32'H7146: READ <= 8'Hd7;
      32'H7147: READ <= 8'Hd7;
      32'H7148: READ <= 8'Hd6;
      32'H7149: READ <= 8'Hd5;
      32'H7150: READ <= 8'Hd2;
      32'H7151: READ <= 8'Hd1;
      32'H7152: READ <= 8'Hcf;
      32'H7153: READ <= 8'Hd1;
      32'H7154: READ <= 8'Hd6;
      32'H7155: READ <= 8'Hd8;
      32'H7156: READ <= 8'Hd7;
      32'H7157: READ <= 8'Hd9;
      32'H7158: READ <= 8'Hd6;
      32'H7159: READ <= 8'Hd1;
      32'H7160: READ <= 8'Hcd;
      32'H7161: READ <= 8'Hc6;
      32'H7162: READ <= 8'Hbe;
      32'H7163: READ <= 8'Hb1;
      32'H7164: READ <= 8'Ha4;
      32'H7165: READ <= 8'H9b;
      32'H7166: READ <= 8'H93;
      32'H7167: READ <= 8'H8c;
      32'H7168: READ <= 8'H88;
      32'H7169: READ <= 8'H85;
      32'H7170: READ <= 8'H80;
      32'H7171: READ <= 8'H7b;
      32'H7172: READ <= 8'H7a;
      32'H7173: READ <= 8'H77;
      32'H7174: READ <= 8'H75;
      32'H7175: READ <= 8'H75;
      32'H7176: READ <= 8'H75;
      32'H7177: READ <= 8'H76;
      32'H7178: READ <= 8'H77;
      32'H7179: READ <= 8'H78;
      32'H7180: READ <= 8'H79;
      32'H7181: READ <= 8'H7a;
      32'H7182: READ <= 8'H7b;
      32'H7183: READ <= 8'H7b;
      32'H7184: READ <= 8'H7d;
      32'H7185: READ <= 8'H7d;
      32'H7186: READ <= 8'H7e;
      32'H7187: READ <= 8'H80;
      32'H7188: READ <= 8'H7f;
      32'H7189: READ <= 8'H81;
      32'H7190: READ <= 8'H82;
      32'H7191: READ <= 8'H82;
      32'H7192: READ <= 8'H82;
      32'H7193: READ <= 8'H84;
      32'H7194: READ <= 8'H85;
      32'H7195: READ <= 8'H86;
      32'H7196: READ <= 8'H86;
      32'H7197: READ <= 8'H86;
      32'H7198: READ <= 8'H87;
      32'H7199: READ <= 8'H87;
      32'H7200: READ <= 8'H75;
      32'H7201: READ <= 8'H76;
      32'H7202: READ <= 8'H76;
      32'H7203: READ <= 8'H75;
      32'H7204: READ <= 8'H75;
      32'H7205: READ <= 8'H75;
      32'H7206: READ <= 8'H74;
      32'H7207: READ <= 8'H75;
      32'H7208: READ <= 8'H75;
      32'H7209: READ <= 8'H74;
      32'H7210: READ <= 8'H73;
      32'H7211: READ <= 8'H73;
      32'H7212: READ <= 8'H72;
      32'H7213: READ <= 8'H71;
      32'H7214: READ <= 8'H71;
      32'H7215: READ <= 8'H71;
      32'H7216: READ <= 8'H70;
      32'H7217: READ <= 8'H70;
      32'H7218: READ <= 8'H6f;
      32'H7219: READ <= 8'H70;
      32'H7220: READ <= 8'H6f;
      32'H7221: READ <= 8'H6f;
      32'H7222: READ <= 8'H6f;
      32'H7223: READ <= 8'H70;
      32'H7224: READ <= 8'H71;
      32'H7225: READ <= 8'H77;
      32'H7226: READ <= 8'H7e;
      32'H7227: READ <= 8'H86;
      32'H7228: READ <= 8'H8f;
      32'H7229: READ <= 8'H97;
      32'H7230: READ <= 8'H9f;
      32'H7231: READ <= 8'Ha5;
      32'H7232: READ <= 8'Hca;
      32'H7233: READ <= 8'Hbd;
      32'H7234: READ <= 8'Hb2;
      32'H7235: READ <= 8'Hb7;
      32'H7236: READ <= 8'Hc3;
      32'H7237: READ <= 8'Hd0;
      32'H7238: READ <= 8'Hd7;
      32'H7239: READ <= 8'Hda;
      32'H7240: READ <= 8'Hdc;
      32'H7241: READ <= 8'Hdd;
      32'H7242: READ <= 8'Hde;
      32'H7243: READ <= 8'Hdb;
      32'H7244: READ <= 8'Hd9;
      32'H7245: READ <= 8'Hd8;
      32'H7246: READ <= 8'Hd9;
      32'H7247: READ <= 8'Hd9;
      32'H7248: READ <= 8'Hd9;
      32'H7249: READ <= 8'Hd8;
      32'H7250: READ <= 8'Hd7;
      32'H7251: READ <= 8'Hd6;
      32'H7252: READ <= 8'Hd6;
      32'H7253: READ <= 8'Hda;
      32'H7254: READ <= 8'Hdb;
      32'H7255: READ <= 8'Hdd;
      32'H7256: READ <= 8'Hde;
      32'H7257: READ <= 8'Hdb;
      32'H7258: READ <= 8'Hd7;
      32'H7259: READ <= 8'Hd3;
      32'H7260: READ <= 8'Hcf;
      32'H7261: READ <= 8'Hc9;
      32'H7262: READ <= 8'Hc0;
      32'H7263: READ <= 8'Hb5;
      32'H7264: READ <= 8'Ha9;
      32'H7265: READ <= 8'H9d;
      32'H7266: READ <= 8'H96;
      32'H7267: READ <= 8'H90;
      32'H7268: READ <= 8'H8b;
      32'H7269: READ <= 8'H87;
      32'H7270: READ <= 8'H83;
      32'H7271: READ <= 8'H7e;
      32'H7272: READ <= 8'H7b;
      32'H7273: READ <= 8'H78;
      32'H7274: READ <= 8'H76;
      32'H7275: READ <= 8'H76;
      32'H7276: READ <= 8'H75;
      32'H7277: READ <= 8'H75;
      32'H7278: READ <= 8'H77;
      32'H7279: READ <= 8'H78;
      32'H7280: READ <= 8'H78;
      32'H7281: READ <= 8'H79;
      32'H7282: READ <= 8'H7b;
      32'H7283: READ <= 8'H7b;
      32'H7284: READ <= 8'H7c;
      32'H7285: READ <= 8'H7c;
      32'H7286: READ <= 8'H7e;
      32'H7287: READ <= 8'H7f;
      32'H7288: READ <= 8'H80;
      32'H7289: READ <= 8'H81;
      32'H7290: READ <= 8'H82;
      32'H7291: READ <= 8'H82;
      32'H7292: READ <= 8'H83;
      32'H7293: READ <= 8'H84;
      32'H7294: READ <= 8'H85;
      32'H7295: READ <= 8'H85;
      32'H7296: READ <= 8'H85;
      32'H7297: READ <= 8'H86;
      32'H7298: READ <= 8'H87;
      32'H7299: READ <= 8'H87;
      32'H7300: READ <= 8'H76;
      32'H7301: READ <= 8'H76;
      32'H7302: READ <= 8'H76;
      32'H7303: READ <= 8'H76;
      32'H7304: READ <= 8'H76;
      32'H7305: READ <= 8'H76;
      32'H7306: READ <= 8'H75;
      32'H7307: READ <= 8'H75;
      32'H7308: READ <= 8'H75;
      32'H7309: READ <= 8'H74;
      32'H7310: READ <= 8'H74;
      32'H7311: READ <= 8'H74;
      32'H7312: READ <= 8'H73;
      32'H7313: READ <= 8'H72;
      32'H7314: READ <= 8'H73;
      32'H7315: READ <= 8'H71;
      32'H7316: READ <= 8'H71;
      32'H7317: READ <= 8'H70;
      32'H7318: READ <= 8'H70;
      32'H7319: READ <= 8'H70;
      32'H7320: READ <= 8'H70;
      32'H7321: READ <= 8'H70;
      32'H7322: READ <= 8'H70;
      32'H7323: READ <= 8'H70;
      32'H7324: READ <= 8'H72;
      32'H7325: READ <= 8'H77;
      32'H7326: READ <= 8'H7f;
      32'H7327: READ <= 8'H88;
      32'H7328: READ <= 8'H90;
      32'H7329: READ <= 8'H99;
      32'H7330: READ <= 8'Ha1;
      32'H7331: READ <= 8'Had;
      32'H7332: READ <= 8'Hd0;
      32'H7333: READ <= 8'Hb5;
      32'H7334: READ <= 8'Ha0;
      32'H7335: READ <= 8'Hb4;
      32'H7336: READ <= 8'Hb6;
      32'H7337: READ <= 8'Hc8;
      32'H7338: READ <= 8'Hd3;
      32'H7339: READ <= 8'Hd9;
      32'H7340: READ <= 8'Hdb;
      32'H7341: READ <= 8'Hdc;
      32'H7342: READ <= 8'Hde;
      32'H7343: READ <= 8'Hdd;
      32'H7344: READ <= 8'Hdc;
      32'H7345: READ <= 8'Hdc;
      32'H7346: READ <= 8'Hdd;
      32'H7347: READ <= 8'Hdd;
      32'H7348: READ <= 8'Hdb;
      32'H7349: READ <= 8'Hdb;
      32'H7350: READ <= 8'Hdb;
      32'H7351: READ <= 8'Hdc;
      32'H7352: READ <= 8'Hdc;
      32'H7353: READ <= 8'Hde;
      32'H7354: READ <= 8'Hde;
      32'H7355: READ <= 8'Hdf;
      32'H7356: READ <= 8'He0;
      32'H7357: READ <= 8'Hdd;
      32'H7358: READ <= 8'Hd9;
      32'H7359: READ <= 8'Hd5;
      32'H7360: READ <= 8'Hd0;
      32'H7361: READ <= 8'Hcc;
      32'H7362: READ <= 8'Hc4;
      32'H7363: READ <= 8'Hb9;
      32'H7364: READ <= 8'Hac;
      32'H7365: READ <= 8'Ha1;
      32'H7366: READ <= 8'H99;
      32'H7367: READ <= 8'H92;
      32'H7368: READ <= 8'H8e;
      32'H7369: READ <= 8'H89;
      32'H7370: READ <= 8'H85;
      32'H7371: READ <= 8'H80;
      32'H7372: READ <= 8'H7d;
      32'H7373: READ <= 8'H7a;
      32'H7374: READ <= 8'H77;
      32'H7375: READ <= 8'H78;
      32'H7376: READ <= 8'H76;
      32'H7377: READ <= 8'H76;
      32'H7378: READ <= 8'H77;
      32'H7379: READ <= 8'H78;
      32'H7380: READ <= 8'H79;
      32'H7381: READ <= 8'H79;
      32'H7382: READ <= 8'H7b;
      32'H7383: READ <= 8'H7b;
      32'H7384: READ <= 8'H7c;
      32'H7385: READ <= 8'H7d;
      32'H7386: READ <= 8'H7e;
      32'H7387: READ <= 8'H7e;
      32'H7388: READ <= 8'H80;
      32'H7389: READ <= 8'H80;
      32'H7390: READ <= 8'H81;
      32'H7391: READ <= 8'H83;
      32'H7392: READ <= 8'H83;
      32'H7393: READ <= 8'H83;
      32'H7394: READ <= 8'H85;
      32'H7395: READ <= 8'H85;
      32'H7396: READ <= 8'H86;
      32'H7397: READ <= 8'H86;
      32'H7398: READ <= 8'H87;
      32'H7399: READ <= 8'H86;
      32'H7400: READ <= 8'H76;
      32'H7401: READ <= 8'H76;
      32'H7402: READ <= 8'H76;
      32'H7403: READ <= 8'H75;
      32'H7404: READ <= 8'H76;
      32'H7405: READ <= 8'H76;
      32'H7406: READ <= 8'H76;
      32'H7407: READ <= 8'H75;
      32'H7408: READ <= 8'H76;
      32'H7409: READ <= 8'H75;
      32'H7410: READ <= 8'H74;
      32'H7411: READ <= 8'H74;
      32'H7412: READ <= 8'H74;
      32'H7413: READ <= 8'H73;
      32'H7414: READ <= 8'H73;
      32'H7415: READ <= 8'H71;
      32'H7416: READ <= 8'H71;
      32'H7417: READ <= 8'H71;
      32'H7418: READ <= 8'H70;
      32'H7419: READ <= 8'H70;
      32'H7420: READ <= 8'H70;
      32'H7421: READ <= 8'H70;
      32'H7422: READ <= 8'H70;
      32'H7423: READ <= 8'H71;
      32'H7424: READ <= 8'H74;
      32'H7425: READ <= 8'H78;
      32'H7426: READ <= 8'H7f;
      32'H7427: READ <= 8'H88;
      32'H7428: READ <= 8'H91;
      32'H7429: READ <= 8'H9b;
      32'H7430: READ <= 8'Ha3;
      32'H7431: READ <= 8'Hb6;
      32'H7432: READ <= 8'Hcd;
      32'H7433: READ <= 8'Hb5;
      32'H7434: READ <= 8'H9c;
      32'H7435: READ <= 8'Hab;
      32'H7436: READ <= 8'Hb6;
      32'H7437: READ <= 8'Hc3;
      32'H7438: READ <= 8'Hce;
      32'H7439: READ <= 8'Hd7;
      32'H7440: READ <= 8'Hda;
      32'H7441: READ <= 8'Hdc;
      32'H7442: READ <= 8'Hde;
      32'H7443: READ <= 8'Hdd;
      32'H7444: READ <= 8'Hdc;
      32'H7445: READ <= 8'Hdd;
      32'H7446: READ <= 8'Hde;
      32'H7447: READ <= 8'Hdf;
      32'H7448: READ <= 8'Hde;
      32'H7449: READ <= 8'Hde;
      32'H7450: READ <= 8'Hde;
      32'H7451: READ <= 8'Hdf;
      32'H7452: READ <= 8'Hdf;
      32'H7453: READ <= 8'He0;
      32'H7454: READ <= 8'He1;
      32'H7455: READ <= 8'He2;
      32'H7456: READ <= 8'He1;
      32'H7457: READ <= 8'Hde;
      32'H7458: READ <= 8'Hdb;
      32'H7459: READ <= 8'Hd6;
      32'H7460: READ <= 8'Hd2;
      32'H7461: READ <= 8'Hcd;
      32'H7462: READ <= 8'Hc6;
      32'H7463: READ <= 8'Hbb;
      32'H7464: READ <= 8'Hb0;
      32'H7465: READ <= 8'Ha4;
      32'H7466: READ <= 8'H9b;
      32'H7467: READ <= 8'H93;
      32'H7468: READ <= 8'H8f;
      32'H7469: READ <= 8'H8b;
      32'H7470: READ <= 8'H87;
      32'H7471: READ <= 8'H82;
      32'H7472: READ <= 8'H7f;
      32'H7473: READ <= 8'H7d;
      32'H7474: READ <= 8'H7a;
      32'H7475: READ <= 8'H77;
      32'H7476: READ <= 8'H76;
      32'H7477: READ <= 8'H77;
      32'H7478: READ <= 8'H77;
      32'H7479: READ <= 8'H77;
      32'H7480: READ <= 8'H78;
      32'H7481: READ <= 8'H79;
      32'H7482: READ <= 8'H7b;
      32'H7483: READ <= 8'H7c;
      32'H7484: READ <= 8'H7c;
      32'H7485: READ <= 8'H7d;
      32'H7486: READ <= 8'H7e;
      32'H7487: READ <= 8'H7e;
      32'H7488: READ <= 8'H7f;
      32'H7489: READ <= 8'H81;
      32'H7490: READ <= 8'H81;
      32'H7491: READ <= 8'H82;
      32'H7492: READ <= 8'H83;
      32'H7493: READ <= 8'H83;
      32'H7494: READ <= 8'H85;
      32'H7495: READ <= 8'H85;
      32'H7496: READ <= 8'H85;
      32'H7497: READ <= 8'H86;
      32'H7498: READ <= 8'H86;
      32'H7499: READ <= 8'H86;
      default: READ <= 8'bx;
  endcase
end

endmodule
